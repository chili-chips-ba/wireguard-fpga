-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 984
entity tb_0CLK_3cb1e4cb is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 global_to_module : in tb_global_to_module_t;
 module_to_global : out tb_module_to_global_t;
 return_output : out axis128_t_stream_t);
end tb_0CLK_3cb1e4cb;
architecture arch of tb_0CLK_3cb1e4cb is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal input_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal ciphertext_in_stream : uint8_t_144 := (others => to_unsigned(0, 8));
signal ciphertext_remaining_in : unsigned(31 downto 0) := to_unsigned(0, 32);
signal cycle_counter : unsigned(31 downto 0) := to_unsigned(0, 32);
signal output_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_size : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_remaining_out : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_expected : uint8_t_128 := (others => to_unsigned(0, 8));
signal tag_match_checked : unsigned(0 downto 0) := to_unsigned(0, 1);
signal chacha20poly1305_decrypt_axis_in : axis128_t_stream_t := axis128_t_stream_t_NULL;
signal REG_COMB_input_packet_count : unsigned(31 downto 0);
signal REG_COMB_ciphertext_in_stream : uint8_t_144;
signal REG_COMB_ciphertext_remaining_in : unsigned(31 downto 0);
signal REG_COMB_cycle_counter : unsigned(31 downto 0);
signal REG_COMB_output_packet_count : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_size : unsigned(31 downto 0);
signal REG_COMB_plaintext_remaining_out : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_expected : uint8_t_128;
signal REG_COMB_tag_match_checked : unsigned(0 downto 0);
signal REG_COMB_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;

-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l179_c8_09da]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l180_c1_7711]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : uint8_t_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : uint8_t_144;

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165[chacha20poly1305_decrypt_tb_c_l181_c9_9165]
signal printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165_CLOCK_ENABLE : unsigned(0 downto 0);

-- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l183_c117_2a9b]
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_x : unsigned(255 downto 0);
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output : unsigned(255 downto 0);

-- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l183_c148_c11e]
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_x : unsigned(255 downto 0);
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output : unsigned(255 downto 0);

-- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l183_c179_093b]
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_x : unsigned(255 downto 0);
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output : unsigned(255 downto 0);

-- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l183_c210_a1cc]
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_x : unsigned(255 downto 0);
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output : unsigned(255 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l183_c241_1fac]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_x : unsigned(255 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output : unsigned(255 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l183_c272_c1b2]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_x : unsigned(255 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output : unsigned(255 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l183_c302_1489]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_x : unsigned(255 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output : unsigned(255 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l183_c332_d4d8]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_x : unsigned(255 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output : unsigned(255 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743[chacha20poly1305_decrypt_tb_c_l183_c64_5743]
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg3 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg4 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg5 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg6 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg7 : unsigned(31 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l184_c100_1c53]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_x : unsigned(95 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output : unsigned(95 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l184_c130_4c71]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_x : unsigned(95 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output : unsigned(95 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l184_c160_32aa]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_x : unsigned(95 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output : unsigned(95 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1[chacha20poly1305_decrypt_tb_c_l184_c65_d1b1]
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg2 : unsigned(31 downto 0);

-- print_aad[chacha20poly1305_decrypt_tb_c_l185_c9_3334]
signal print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_CLOCK_ENABLE : unsigned(0 downto 0);
signal print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad : uint8_t_32;
signal print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad_len : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l189_c32_0b54]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l190_c35_6769]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0[chacha20poly1305_decrypt_tb_c_l191_c9_8ae0]
signal printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg1 : unsigned(31 downto 0);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l194_c30_26c6]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l198_c34_97d4]
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_0 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_1 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output : uint8_t_array_128_t;

-- printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0[chacha20poly1305_decrypt_tb_c_l200_c9_53d0]
signal printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l205_c9_1d2f]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_right : unsigned(0 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output : unsigned(0 downto 0);

-- BIN_OP_MOD[chacha20poly1305_decrypt_tb_c_l205_c31_26fa]
signal BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_left : unsigned(31 downto 0);
signal BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_right : unsigned(4 downto 0);
signal BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output : unsigned(4 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l205_c31_15f7]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_left : unsigned(4 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l205_c9_cfd1]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output : unsigned(0 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l205_c59_fd85]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_right : unsigned(0 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l205_c9_2fad]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l205_c1_c273]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68[chacha20poly1305_decrypt_tb_c_l206_c9_6d68]
signal printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l213_c8_7e08]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_right : unsigned(0 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l214_c1_8bf9]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(31 downto 0);

-- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4]
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : axis128_t_stream_t;

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac]
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);

-- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l227_c56_6fd6]
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_left : unsigned(31 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_right : unsigned(4 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l230_c12_c373]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l231_c1_de39]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(31 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l232_c176_e3c5]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l232_c207_f310]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l232_c237_0c4e]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l232_c267_3cbf]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1[chacha20poly1305_decrypt_tb_c_l232_c108_5fc1]
signal printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg3 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l234_c1_b6b6]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output : unsigned(0 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d[chacha20poly1305_decrypt_tb_c_l235_c17_7f1d]
signal printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l237_c17_bf36]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l239_c17_0476]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output : unsigned(31 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l248_c8_f415]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l249_c1_f913]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(31 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l251_c169_6c9e]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l251_c200_2176]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l251_c230_8416]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l251_c260_51b2]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b[chacha20poly1305_decrypt_tb_c_l251_c105_b34b]
signal printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg3 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f]
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l268_c1_2dea]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l275_c1_88c6]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l269_c16_4da1]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_right : unsigned(4 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l269_c1_5c29]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l271_c1_bc29]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l269_c13_ea14]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd[chacha20poly1305_decrypt_tb_c_l270_c17_aafd]
signal printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_CLOCK_ENABLE : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b[chacha20poly1305_decrypt_tb_c_l272_c17_fb9b]
signal printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_arg0 : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l276_c16_9117]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l276_c1_6034]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d[chacha20poly1305_decrypt_tb_c_l277_c18_784d]
signal printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l279_c17_fb4e]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l286_c9_4b3b]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output : unsigned(0 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l286_c41_a2b3]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l286_c9_e09e]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output : unsigned(0 downto 0);

-- UNARY_OP_NOT[chacha20poly1305_decrypt_tb_c_l286_c69_ef49]
signal UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l286_c9_21ab]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l287_c1_acb3]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : uint8_t_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : uint8_t_144;

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);

-- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1]
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l288_c13_fe56]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_left : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l289_c1_ec75]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l291_c1_cbc7]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695[chacha20poly1305_decrypt_tb_c_l290_c13_9695]
signal printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_arg0 : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a[chacha20poly1305_decrypt_tb_c_l292_c13_395a]
signal printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l296_c9_e3e9]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output : unsigned(32 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l297_c12_2242]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l298_c1_84a2]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : uint8_t_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : uint8_t_144;

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l300_c17_b9d8]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_right : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l300_c1_bafe]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output : unsigned(0 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : uint8_t_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : uint8_t_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : uint8_t_144;

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l302_c40_0822]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l303_c43_94e2]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4[chacha20poly1305_decrypt_tb_c_l304_c17_01e4]
signal printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg1 : unsigned(31 downto 0);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l307_c38_317b]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l311_c42_328d]
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_0 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_1 : uint8_t_128;
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output : uint8_t_array_128_t;

-- printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e[chacha20poly1305_decrypt_tb_c_l313_c17_391e]
signal printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l320_c9_eb04]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_right : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output : unsigned(0 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l320_c5_c1e4]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l324_c5_e824]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_right : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint8_t_144_uint8_t_144_a26f( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_b938( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;
      base(80) := ref_toks_81;
      base(81) := ref_toks_82;
      base(82) := ref_toks_83;
      base(83) := ref_toks_84;
      base(84) := ref_toks_85;
      base(85) := ref_toks_86;
      base(86) := ref_toks_87;
      base(87) := ref_toks_88;
      base(88) := ref_toks_89;
      base(89) := ref_toks_90;
      base(90) := ref_toks_91;
      base(91) := ref_toks_92;
      base(92) := ref_toks_93;
      base(93) := ref_toks_94;
      base(94) := ref_toks_95;
      base(95) := ref_toks_96;

      return_output := base;
      return return_output; 
end function;

function uint8_array32_be( x : uint8_t_32) return unsigned is

  --variable x : uint8_t_32;
  variable return_output : unsigned(255 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15)&x(16)&x(17)&x(18)&x(19)&x(20)&x(21)&x(22)&x(23)&x(24)&x(25)&x(26)&x(27)&x(28)&x(29)&x(30)&x(31);
return return_output;
end function;

function uint8_array12_be( x : uint8_t_12) return unsigned is

  --variable x : uint8_t_12;
  variable return_output : unsigned(95 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11);
return return_output;
end function;

function CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_16 is
 
  variable base : axis128_t_stream_t; 
  variable return_output : uint8_t_16;
begin
      base.data.tdata(0) := ref_toks_0;
      base.data.tdata(1) := ref_toks_1;
      base.data.tdata(2) := ref_toks_2;
      base.data.tdata(3) := ref_toks_3;
      base.data.tdata(4) := ref_toks_4;
      base.data.tdata(5) := ref_toks_5;
      base.data.tdata(6) := ref_toks_6;
      base.data.tdata(7) := ref_toks_7;
      base.data.tdata(8) := ref_toks_8;
      base.data.tdata(9) := ref_toks_9;
      base.data.tdata(10) := ref_toks_10;
      base.data.tdata(11) := ref_toks_11;
      base.data.tdata(12) := ref_toks_12;
      base.data.tdata(13) := ref_toks_13;
      base.data.tdata(14) := ref_toks_14;
      base.data.tdata(15) := ref_toks_15;

      return_output := base.data.tdata;
      return return_output; 
end function;

function uint8_array16_be( x : uint8_t_16) return unsigned is

  --variable x : uint8_t_16;
  variable return_output : unsigned(127 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15);
return return_output;
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base.data.tkeep(0) := ref_toks_0;
      base.data.tdata(0) := ref_toks_1;
      base.data.tkeep(1) := ref_toks_2;
      base.data.tdata(1) := ref_toks_3;
      base.data.tkeep(2) := ref_toks_4;
      base.data.tdata(2) := ref_toks_5;
      base.data.tkeep(3) := ref_toks_6;
      base.data.tdata(3) := ref_toks_7;
      base.data.tkeep(4) := ref_toks_8;
      base.data.tdata(4) := ref_toks_9;
      base.data.tkeep(5) := ref_toks_10;
      base.data.tdata(5) := ref_toks_11;
      base.data.tkeep(6) := ref_toks_12;
      base.data.tdata(6) := ref_toks_13;
      base.data.tkeep(7) := ref_toks_14;
      base.data.tdata(7) := ref_toks_15;
      base.data.tkeep(8) := ref_toks_16;
      base.data.tdata(8) := ref_toks_17;
      base.data.tkeep(9) := ref_toks_18;
      base.data.tdata(9) := ref_toks_19;
      base.data.tkeep(10) := ref_toks_20;
      base.data.tdata(10) := ref_toks_21;
      base.data.tkeep(11) := ref_toks_22;
      base.data.tdata(11) := ref_toks_23;
      base.data.tkeep(12) := ref_toks_24;
      base.data.tdata(12) := ref_toks_25;
      base.data.tkeep(13) := ref_toks_26;
      base.data.tdata(13) := ref_toks_27;
      base.data.tkeep(14) := ref_toks_28;
      base.data.tdata(14) := ref_toks_29;
      base.data.tkeep(15) := ref_toks_30;
      base.data.tdata(15) := ref_toks_31;
      base.data.tlast := ref_toks_32;
      base.valid := ref_toks_33;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee( ref_toks_0 : axis128_t_stream_t;
 ref_toks_1 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base := ref_toks_0;
      base.valid := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_32_uint8_t_32_1367( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned) return uint8_t_32 is
 
  variable base : uint8_t_32; 
  variable return_output : uint8_t_32;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;
      base(12) := ref_toks_12;
      base(13) := ref_toks_13;
      base(14) := ref_toks_14;
      base(15) := ref_toks_15;
      base(16) := ref_toks_16;
      base(17) := ref_toks_17;
      base(18) := ref_toks_18;
      base(19) := ref_toks_19;
      base(20) := ref_toks_20;
      base(21) := ref_toks_21;
      base(22) := ref_toks_22;
      base(23) := ref_toks_23;
      base(24) := ref_toks_24;
      base(25) := ref_toks_25;
      base(26) := ref_toks_26;
      base(27) := ref_toks_27;
      base(28) := ref_toks_28;
      base(29) := ref_toks_29;
      base(30) := ref_toks_30;
      base(31) := ref_toks_31;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return uint8_t_12 is
 
  variable base : uint8_t_12; 
  variable return_output : uint8_t_12;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_128_uint8_t_128_7166( ref_toks_0 : uint8_t_128;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned) return uint8_t_128 is
 
  variable base : uint8_t_128; 
  variable return_output : uint8_t_128;
begin
      base := ref_toks_0;
      base(103) := ref_toks_1;
      base(48) := ref_toks_2;
      base(57) := ref_toks_3;
      base(54) := ref_toks_4;
      base(63) := ref_toks_5;
      base(8) := ref_toks_6;
      base(72) := ref_toks_7;
      base(17) := ref_toks_8;
      base(81) := ref_toks_9;
      base(26) := ref_toks_10;
      base(23) := ref_toks_11;
      base(90) := ref_toks_12;
      base(87) := ref_toks_13;
      base(32) := ref_toks_14;
      base(96) := ref_toks_15;
      base(41) := ref_toks_16;
      base(105) := ref_toks_17;
      base(50) := ref_toks_18;
      base(47) := ref_toks_19;
      base(59) := ref_toks_20;
      base(111) := ref_toks_21;
      base(56) := ref_toks_22;
      base(1) := ref_toks_23;
      base(65) := ref_toks_24;
      base(10) := ref_toks_25;
      base(74) := ref_toks_26;
      base(19) := ref_toks_27;
      base(16) := ref_toks_28;
      base(83) := ref_toks_29;
      base(80) := ref_toks_30;
      base(25) := ref_toks_31;
      base(89) := ref_toks_32;
      base(34) := ref_toks_33;
      base(98) := ref_toks_34;
      base(43) := ref_toks_35;
      base(107) := ref_toks_36;
      base(52) := ref_toks_37;
      base(49) := ref_toks_38;
      base(58) := ref_toks_39;
      base(3) := ref_toks_40;
      base(67) := ref_toks_41;
      base(12) := ref_toks_42;
      base(9) := ref_toks_43;
      base(76) := ref_toks_44;
      base(73) := ref_toks_45;
      base(18) := ref_toks_46;
      base(85) := ref_toks_47;
      base(82) := ref_toks_48;
      base(27) := ref_toks_49;
      base(91) := ref_toks_50;
      base(36) := ref_toks_51;
      base(100) := ref_toks_52;
      base(45) := ref_toks_53;
      base(30) := ref_toks_54;
      base(109) := ref_toks_55;
      base(42) := ref_toks_56;
      base(106) := ref_toks_57;
      base(51) := ref_toks_58;
      base(60) := ref_toks_59;
      base(5) := ref_toks_60;
      base(2) := ref_toks_61;
      base(69) := ref_toks_62;
      base(14) := ref_toks_63;
      base(66) := ref_toks_64;
      base(11) := ref_toks_65;
      base(78) := ref_toks_66;
      base(75) := ref_toks_67;
      base(20) := ref_toks_68;
      base(84) := ref_toks_69;
      base(29) := ref_toks_70;
      base(93) := ref_toks_71;
      base(38) := ref_toks_72;
      base(102) := ref_toks_73;
      base(35) := ref_toks_74;
      base(99) := ref_toks_75;
      base(44) := ref_toks_76;
      base(108) := ref_toks_77;
      base(53) := ref_toks_78;
      base(62) := ref_toks_79;
      base(7) := ref_toks_80;
      base(4) := ref_toks_81;
      base(71) := ref_toks_82;
      base(68) := ref_toks_83;
      base(13) := ref_toks_84;
      base(77) := ref_toks_85;
      base(22) := ref_toks_86;
      base(86) := ref_toks_87;
      base(31) := ref_toks_88;
      base(95) := ref_toks_89;
      base(28) := ref_toks_90;
      base(40) := ref_toks_91;
      base(92) := ref_toks_92;
      base(104) := ref_toks_93;
      base(37) := ref_toks_94;
      base(101) := ref_toks_95;
      base(46) := ref_toks_96;
      base(110) := ref_toks_97;
      base(55) := ref_toks_98;
      base(0) := ref_toks_99;
      base(64) := ref_toks_100;
      base(61) := ref_toks_101;
      base(6) := ref_toks_102;
      base(70) := ref_toks_103;
      base(15) := ref_toks_104;
      base(79) := ref_toks_105;
      base(24) := ref_toks_106;
      base(88) := ref_toks_107;
      base(21) := ref_toks_108;
      base(33) := ref_toks_109;
      base(97) := ref_toks_110;
      base(94) := ref_toks_111;
      base(39) := ref_toks_112;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned;
 ref_toks_113 : unsigned;
 ref_toks_114 : unsigned;
 ref_toks_115 : unsigned;
 ref_toks_116 : unsigned;
 ref_toks_117 : unsigned;
 ref_toks_118 : unsigned;
 ref_toks_119 : unsigned;
 ref_toks_120 : unsigned;
 ref_toks_121 : unsigned;
 ref_toks_122 : unsigned;
 ref_toks_123 : unsigned;
 ref_toks_124 : unsigned;
 ref_toks_125 : unsigned;
 ref_toks_126 : unsigned;
 ref_toks_127 : unsigned;
 ref_toks_128 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(113) := ref_toks_1;
      base(122) := ref_toks_2;
      base(15) := ref_toks_3;
      base(79) := ref_toks_4;
      base(24) := ref_toks_5;
      base(88) := ref_toks_6;
      base(33) := ref_toks_7;
      base(97) := ref_toks_8;
      base(42) := ref_toks_9;
      base(106) := ref_toks_10;
      base(51) := ref_toks_11;
      base(115) := ref_toks_12;
      base(8) := ref_toks_13;
      base(72) := ref_toks_14;
      base(17) := ref_toks_15;
      base(81) := ref_toks_16;
      base(26) := ref_toks_17;
      base(90) := ref_toks_18;
      base(35) := ref_toks_19;
      base(99) := ref_toks_20;
      base(44) := ref_toks_21;
      base(108) := ref_toks_22;
      base(1) := ref_toks_23;
      base(65) := ref_toks_24;
      base(10) := ref_toks_25;
      base(74) := ref_toks_26;
      base(19) := ref_toks_27;
      base(83) := ref_toks_28;
      base(28) := ref_toks_29;
      base(92) := ref_toks_30;
      base(37) := ref_toks_31;
      base(101) := ref_toks_32;
      base(58) := ref_toks_33;
      base(3) := ref_toks_34;
      base(67) := ref_toks_35;
      base(12) := ref_toks_36;
      base(76) := ref_toks_37;
      base(21) := ref_toks_38;
      base(85) := ref_toks_39;
      base(30) := ref_toks_40;
      base(94) := ref_toks_41;
      base(60) := ref_toks_42;
      base(5) := ref_toks_43;
      base(124) := ref_toks_44;
      base(69) := ref_toks_45;
      base(14) := ref_toks_46;
      base(78) := ref_toks_47;
      base(23) := ref_toks_48;
      base(87) := ref_toks_49;
      base(32) := ref_toks_50;
      base(96) := ref_toks_51;
      base(53) := ref_toks_52;
      base(117) := ref_toks_53;
      base(62) := ref_toks_54;
      base(7) := ref_toks_55;
      base(126) := ref_toks_56;
      base(71) := ref_toks_57;
      base(16) := ref_toks_58;
      base(80) := ref_toks_59;
      base(25) := ref_toks_60;
      base(89) := ref_toks_61;
      base(46) := ref_toks_62;
      base(110) := ref_toks_63;
      base(55) := ref_toks_64;
      base(0) := ref_toks_65;
      base(119) := ref_toks_66;
      base(64) := ref_toks_67;
      base(9) := ref_toks_68;
      base(73) := ref_toks_69;
      base(18) := ref_toks_70;
      base(82) := ref_toks_71;
      base(39) := ref_toks_72;
      base(103) := ref_toks_73;
      base(48) := ref_toks_74;
      base(112) := ref_toks_75;
      base(57) := ref_toks_76;
      base(2) := ref_toks_77;
      base(121) := ref_toks_78;
      base(66) := ref_toks_79;
      base(11) := ref_toks_80;
      base(75) := ref_toks_81;
      base(41) := ref_toks_82;
      base(105) := ref_toks_83;
      base(50) := ref_toks_84;
      base(114) := ref_toks_85;
      base(59) := ref_toks_86;
      base(4) := ref_toks_87;
      base(123) := ref_toks_88;
      base(68) := ref_toks_89;
      base(77) := ref_toks_90;
      base(34) := ref_toks_91;
      base(98) := ref_toks_92;
      base(43) := ref_toks_93;
      base(107) := ref_toks_94;
      base(52) := ref_toks_95;
      base(116) := ref_toks_96;
      base(61) := ref_toks_97;
      base(6) := ref_toks_98;
      base(125) := ref_toks_99;
      base(70) := ref_toks_100;
      base(27) := ref_toks_101;
      base(91) := ref_toks_102;
      base(36) := ref_toks_103;
      base(100) := ref_toks_104;
      base(45) := ref_toks_105;
      base(109) := ref_toks_106;
      base(54) := ref_toks_107;
      base(118) := ref_toks_108;
      base(63) := ref_toks_109;
      base(127) := ref_toks_110;
      base(20) := ref_toks_111;
      base(84) := ref_toks_112;
      base(29) := ref_toks_113;
      base(93) := ref_toks_114;
      base(38) := ref_toks_115;
      base(102) := ref_toks_116;
      base(47) := ref_toks_117;
      base(111) := ref_toks_118;
      base(56) := ref_toks_119;
      base(120) := ref_toks_120;
      base(13) := ref_toks_121;
      base(22) := ref_toks_122;
      base(86) := ref_toks_123;
      base(31) := ref_toks_124;
      base(95) := ref_toks_125;
      base(40) := ref_toks_126;
      base(104) := ref_toks_127;
      base(49) := ref_toks_128;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165 : entity work.printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165_CLOCK_ENABLE);

-- CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b : 0 clocks latency
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b : entity work.CONST_SR_224_uint256_t_0CLK_de264c78 port map (
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_x,
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output);

-- CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e : 0 clocks latency
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e : entity work.CONST_SR_192_uint256_t_0CLK_de264c78 port map (
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_x,
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output);

-- CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b : 0 clocks latency
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b : entity work.CONST_SR_160_uint256_t_0CLK_de264c78 port map (
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_x,
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output);

-- CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc : 0 clocks latency
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc : entity work.CONST_SR_128_uint256_t_0CLK_de264c78 port map (
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_x,
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac : entity work.CONST_SR_96_uint256_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2 : entity work.CONST_SR_64_uint256_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489 : entity work.CONST_SR_32_uint256_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8 : entity work.CONST_SR_0_uint256_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743 : entity work.printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg0,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg1,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg2,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg3,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg4,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg5,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg6,
printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg7);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53 : entity work.CONST_SR_64_uint96_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71 : entity work.CONST_SR_32_uint96_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa : entity work.CONST_SR_0_uint96_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1 : entity work.printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg0,
printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg1,
printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg2);

-- print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334 : 0 clocks latency
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334 : entity work.print_aad_0CLK_fa355561 port map (
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_CLOCK_ENABLE,
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad,
print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad_len);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54 : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54 : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0 : entity work.printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg0,
printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg1);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4 : 0 clocks latency
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4 : entity work.VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_1,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_var_dim_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0 : entity work.printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg0,
printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f : entity work.BIN_OP_GT_uint32_t_uint1_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output);

-- BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa : 0 clocks latency
BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa : entity work.BIN_OP_MOD_uint32_t_uint5_t_0CLK_29b254e4 port map (
BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_left,
BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_right,
BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7 : entity work.BIN_OP_EQ_uint5_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85 : entity work.BIN_OP_GT_uint32_t_uint1_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68 : entity work.printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg0,
printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08 : entity work.BIN_OP_GT_uint32_t_uint1_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : 0 clocks latency
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4 : entity work.MUX_uint1_t_axis128_t_stream_t_axis128_t_stream_t_0CLK_de264c78 port map (
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

-- BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6 : 0 clocks latency
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6 : entity work.BIN_OP_LTE_uint32_t_uint5_t_0CLK_e595f783 port map (
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_left,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_right,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5 : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5 : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1 : entity work.printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg0,
printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg1,
printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg2,
printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg3);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d : entity work.printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476 : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476 : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416 : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2 : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b : entity work.printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg0,
printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg1,
printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg2,
printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg3);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f : entity work.printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6 : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1 : entity work.BIN_OP_GT_uint32_t_uint5_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29 : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd : entity work.printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_CLOCK_ENABLE);

-- printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b : entity work.printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_arg0);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117 : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d : entity work.printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d_CLOCK_ENABLE);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3 : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3 : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output);

-- UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49 : 0 clocks latency
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_expr,
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : 0 clocks latency
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56 : entity work.BIN_OP_EQ_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7 : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695 : entity work.printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_arg0);

-- printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a : entity work.printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242 : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242 : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8 : entity work.BIN_OP_EQ_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : entity work.MUX_uint1_t_uint8_t_128_uint8_t_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822 : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822 : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4 : entity work.printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg0,
printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg1);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output);

-- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d : 0 clocks latency
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d : entity work.VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_1,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_var_dim_0,
VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e : entity work.printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg0,
printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04 : entity work.BIN_OP_GT_uint32_t_uint32_t_0CLK_380ecc95 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4 : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c : 0 clocks latency
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c : entity work.BIN_OP_MINUS_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_left,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_right,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Registers
 input_packet_count,
 ciphertext_in_stream,
 ciphertext_remaining_in,
 cycle_counter,
 output_packet_count,
 plaintext_out_size,
 plaintext_remaining_out,
 plaintext_out_expected,
 tag_match_checked,
 chacha20poly1305_decrypt_axis_in,
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
 CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output,
 CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output,
 CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output,
 CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output,
 VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output,
 BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
 BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output,
 UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output,
 VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output,
 BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_key : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_nonce : uint8_t_12;
 variable VAR_chacha20poly1305_decrypt_aad : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_aad_len : unsigned(7 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_tags_match : unsigned(0 downto 0);
 variable VAR_key : uint8_t_32;
 variable VAR_nonce : uint8_t_12;
 variable VAR_aad : uint8_t_32;
 variable VAR_aad_len : unsigned(31 downto 0);
 variable VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_fe32_0 : unsigned(31 downto 0);
 variable VAR_plaintexts : uint8_t_2_128;
 variable VAR_plaintext_lens : uint32_t_2;
 variable VAR_input_ciphertext0 : uint8_t_144;
 variable VAR_input_ciphertext1 : uint8_t_144;
 variable VAR_input_ciphertexts : uint8_t_2_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_cf38_return_output : uint8_t_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_fbb8_return_output : uint8_t_144;
 variable VAR_ciphertext_lens : uint32_t_2;
 variable VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l161_c5_13a5 : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l198_c9_532c : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l189_c9_b205 : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_PRINT_32_BYTES_uint : unsigned(255 downto 0);
 variable VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg4 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg5 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg6 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg7 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_x : unsigned(255 downto 0);
 variable VAR_PRINT_12_BYTES_uint : unsigned(95 downto 0);
 variable VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_1caa_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_x : unsigned(95 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad : uint8_t_32;
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad_len : unsigned(31 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output : uint8_t_array_128_t;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_0 : uint8_t_128;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_1 : uint8_t_128;
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output : unsigned(4 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_left : unsigned(4 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iffalse : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond : unsigned(0 downto 0);
 variable VAR_i : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond : unsigned(0 downto 0);
 variable VAR_PRINT_16_BYTES_uint : unsigned(127 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l232_c62_514c_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l232_c45_3245_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_x : unsigned(127 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l237_c17_6bb4 : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output : unsigned(31 downto 0);
 variable VAR_ARRAY_SHIFT_DOWN_i : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l248_c8_c79e_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l251_c58_9d96_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l251_c41_5695_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_x : unsigned(127 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_pos : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_left : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue : unsigned(31 downto 0);
 variable VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55 : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iffalse : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : uint8_t_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l311_c17_860d : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : uint8_t_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l302_c17_010b : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output : uint8_t_array_128_t;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_0 : uint8_t_128;
 variable VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_1 : uint8_t_128;
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_cond : unsigned(0 downto 0);
 variable VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l324_c5_b8b3 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l183_l158_DUPLICATE_0a36_return_output : uint8_t_32;
 variable VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_f336_return_output : uint8_t_12;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_c83e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_37db_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_36c1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_b684_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_efbd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_5abe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_0801_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_eac9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_3f2c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_a48c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_be47_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_ef83_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_671b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_eeb6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_8e59_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_7af8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_7166_chacha20poly1305_decrypt_tb_c_l297_l286_l300_DUPLICATE_f22f_return_output : uint8_t_128;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6_chacha20poly1305_decrypt_tb_c_l286_l300_l297_DUPLICATE_55b0_return_output : uint8_t_144;
 -- State registers comb logic variables
variable REG_VAR_input_packet_count : unsigned(31 downto 0);
variable REG_VAR_ciphertext_in_stream : uint8_t_144;
variable REG_VAR_ciphertext_remaining_in : unsigned(31 downto 0);
variable REG_VAR_cycle_counter : unsigned(31 downto 0);
variable REG_VAR_output_packet_count : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_size : unsigned(31 downto 0);
variable REG_VAR_plaintext_remaining_out : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_expected : uint8_t_128;
variable REG_VAR_tag_match_checked : unsigned(0 downto 0);
variable REG_VAR_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_input_packet_count := input_packet_count;
  REG_VAR_ciphertext_in_stream := ciphertext_in_stream;
  REG_VAR_ciphertext_remaining_in := ciphertext_remaining_in;
  REG_VAR_cycle_counter := cycle_counter;
  REG_VAR_output_packet_count := output_packet_count;
  REG_VAR_plaintext_out_size := plaintext_out_size;
  REG_VAR_plaintext_remaining_out := plaintext_remaining_out;
  REG_VAR_plaintext_out_expected := plaintext_out_expected;
  REG_VAR_tag_match_checked := tag_match_checked;
  REG_VAR_chacha20poly1305_decrypt_axis_in := chacha20poly1305_decrypt_axis_in;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_right := to_unsigned(0, 1);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(12, 32);
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_right := to_unsigned(16, 5);
     VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_right := to_unsigned(20, 5);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_right := to_unsigned(16, 5);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iftrue := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(0, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iffalse := to_unsigned(0, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_0 := to_unsigned(56, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_0 := to_unsigned(56, 32);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(7, 32);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_left := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(1, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(1, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(2, 32);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad := to_byte_array("Additional authenticated data", 32);
     VAR_chacha20poly1305_decrypt_aad := to_byte_array("Additional authenticated data", 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(12, 32);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(15, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(15, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(15, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(1, 32);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_right := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_right := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_right := to_unsigned(1, 1);
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iffalse := to_unsigned(0, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_0 := to_unsigned(80, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_0 := to_unsigned(80, 32);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_right := to_unsigned(16, 5);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_right := to_unsigned(1, 1);
     VAR_chacha20poly1305_decrypt_axis_out_ready := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(2, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iftrue := to_unsigned(0, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_1 := to_unsigned(71, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_1 := to_unsigned(71, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(0, 32);
     VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_fe32_0 := to_unsigned(29, 32);
     VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l161_c5_13a5 := resize(VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_fe32_0, 8);
     VAR_chacha20poly1305_decrypt_aad_len := VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l161_c5_13a5;
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad_len := VAR_aad_len_chacha20poly1305_decrypt_tb_c_l88_c14_fe32_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(4, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(13, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(13, 32);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(9, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(3, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iftrue := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(10, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(11, 32);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_right := to_unsigned(2, 2);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_left := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right := to_signed(14, 32);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_right := to_unsigned(2, 2);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_1 := to_unsigned(96, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_1 := to_unsigned(96, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse := to_unsigned(0, 8);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(14, 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := to_unsigned(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(9, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right := to_signed(4, 32);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_right := to_unsigned(16, 5);
     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l288_c13_fe56] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output;

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_a26f[chacha20poly1305_decrypt_tb_c_l149_c9_cf38] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_cf38_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_a26f(
     (others => to_unsigned(0, 8)),
     to_unsigned(215, 8),
     to_unsigned(30, 8),
     to_unsigned(133, 8),
     to_unsigned(49, 8),
     to_unsigned(110, 8),
     to_unsigned(221, 8),
     to_unsigned(3, 8),
     to_unsigned(242, 8),
     to_unsigned(92, 8),
     to_unsigned(174, 8),
     to_unsigned(198, 8),
     to_unsigned(184, 8),
     to_unsigned(94, 8),
     to_unsigned(232, 8),
     to_unsigned(122, 8),
     to_unsigned(221, 8),
     to_unsigned(225, 8),
     to_unsigned(237, 8),
     to_unsigned(168, 8),
     to_unsigned(104, 8),
     to_unsigned(96, 8),
     to_unsigned(115, 8),
     to_unsigned(11, 8),
     to_unsigned(185, 8),
     to_unsigned(168, 8),
     to_unsigned(235, 8),
     to_unsigned(162, 8),
     to_unsigned(227, 8),
     to_unsigned(117, 8),
     to_unsigned(246, 8),
     to_unsigned(102, 8),
     to_unsigned(196, 8),
     to_unsigned(35, 8),
     to_unsigned(178, 8),
     to_unsigned(235, 8),
     to_unsigned(84, 8),
     to_unsigned(201, 8),
     to_unsigned(250, 8),
     to_unsigned(121, 8),
     to_unsigned(88, 8),
     to_unsigned(152, 8),
     to_unsigned(174, 8),
     to_unsigned(215, 8),
     to_unsigned(124, 8),
     to_unsigned(142, 8),
     to_unsigned(251, 8),
     to_unsigned(38, 8),
     to_unsigned(128, 8),
     to_unsigned(28, 8),
     to_unsigned(119, 8),
     to_unsigned(146, 8),
     to_unsigned(15, 8),
     to_unsigned(219, 8),
     to_unsigned(8, 8),
     to_unsigned(9, 8),
     to_unsigned(110, 8),
     to_unsigned(96, 8),
     to_unsigned(164, 8),
     to_unsigned(133, 8),
     to_unsigned(207, 8),
     to_unsigned(17, 8),
     to_unsigned(184, 8),
     to_unsigned(27, 8),
     to_unsigned(89, 8),
     to_unsigned(93, 8),
     to_unsigned(168, 8),
     to_unsigned(125, 8),
     to_unsigned(106, 8),
     to_unsigned(45, 8),
     to_unsigned(3, 8),
     to_unsigned(201, 8),
     to_unsigned(186, 8),
     to_unsigned(223, 8),
     to_unsigned(92, 8),
     to_unsigned(185, 8),
     to_unsigned(71, 8),
     to_unsigned(116, 8),
     to_unsigned(66, 8),
     to_unsigned(18, 8),
     to_unsigned(63, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_b938[chacha20poly1305_decrypt_tb_c_l150_c9_fbb8] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_fbb8_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_b938(
     (others => to_unsigned(0, 8)),
     to_unsigned(207, 8),
     to_unsigned(18, 8),
     to_unsigned(153, 8),
     to_unsigned(56, 8),
     to_unsigned(109, 8),
     to_unsigned(148, 8),
     to_unsigned(46, 8),
     to_unsigned(223, 8),
     to_unsigned(86, 8),
     to_unsigned(194, 8),
     to_unsigned(230, 8),
     to_unsigned(136, 8),
     to_unsigned(22, 8),
     to_unsigned(245, 8),
     to_unsigned(98, 8),
     to_unsigned(203, 8),
     to_unsigned(225, 8),
     to_unsigned(162, 8),
     to_unsigned(237, 8),
     to_unsigned(76, 8),
     to_unsigned(125, 8),
     to_unsigned(33, 8),
     to_unsigned(38, 8),
     to_unsigned(154, 8),
     to_unsigned(145, 8),
     to_unsigned(170, 8),
     to_unsigned(177, 8),
     to_unsigned(245, 8),
     to_unsigned(58, 8),
     to_unsigned(247, 8),
     to_unsigned(109, 8),
     to_unsigned(193, 8),
     to_unsigned(110, 8),
     to_unsigned(164, 8),
     to_unsigned(226, 8),
     to_unsigned(24, 8),
     to_unsigned(224, 8),
     to_unsigned(235, 8),
     to_unsigned(42, 8),
     to_unsigned(12, 8),
     to_unsigned(203, 8),
     to_unsigned(250, 8),
     to_unsigned(213, 8),
     to_unsigned(96, 8),
     to_unsigned(218, 8),
     to_unsigned(152, 8),
     to_unsigned(26, 8),
     to_unsigned(161, 8),
     to_unsigned(57, 8),
     to_unsigned(77, 8),
     to_unsigned(241, 8),
     to_unsigned(6, 8),
     to_unsigned(215, 8),
     to_unsigned(25, 8),
     to_unsigned(30, 8),
     to_unsigned(111, 8),
     to_unsigned(55, 8),
     to_unsigned(205, 8),
     to_unsigned(247, 8),
     to_unsigned(170, 8),
     to_unsigned(118, 8),
     to_unsigned(205, 8),
     to_unsigned(122, 8),
     to_unsigned(43, 8),
     to_unsigned(152, 8),
     to_unsigned(145, 8),
     to_unsigned(176, 8),
     to_unsigned(58, 8),
     to_unsigned(35, 8),
     to_unsigned(116, 8),
     to_unsigned(207, 8),
     to_unsigned(172, 8),
     to_unsigned(236, 8),
     to_unsigned(106, 8),
     to_unsigned(222, 8),
     to_unsigned(195, 8),
     to_unsigned(78, 8),
     to_unsigned(102, 8),
     to_unsigned(105, 8),
     to_unsigned(120, 8),
     to_unsigned(7, 8),
     to_unsigned(199, 8),
     to_unsigned(227, 8),
     to_unsigned(31, 8),
     to_unsigned(15, 8),
     to_unsigned(235, 8),
     to_unsigned(75, 8),
     to_unsigned(97, 8),
     to_unsigned(234, 8),
     to_unsigned(45, 8),
     to_unsigned(210, 8),
     to_unsigned(164, 8),
     to_unsigned(89, 8),
     to_unsigned(124, 8),
     to_unsigned(174, 8),
     to_unsigned(233, 8));

     -- CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_f336 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_f336_return_output := CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2(
     to_unsigned(7, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(64, 8),
     to_unsigned(65, 8),
     to_unsigned(66, 8),
     to_unsigned(67, 8),
     to_unsigned(68, 8),
     to_unsigned(69, 8),
     to_unsigned(70, 8),
     to_unsigned(71, 8));

     -- CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l183_l158_DUPLICATE_0a36 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l183_l158_DUPLICATE_0a36_return_output := CONST_REF_RD_uint8_t_32_uint8_t_32_1367(
     to_unsigned(128, 8),
     to_unsigned(129, 8),
     to_unsigned(130, 8),
     to_unsigned(131, 8),
     to_unsigned(132, 8),
     to_unsigned(133, 8),
     to_unsigned(134, 8),
     to_unsigned(135, 8),
     to_unsigned(136, 8),
     to_unsigned(137, 8),
     to_unsigned(138, 8),
     to_unsigned(139, 8),
     to_unsigned(140, 8),
     to_unsigned(141, 8),
     to_unsigned(142, 8),
     to_unsigned(143, 8),
     to_unsigned(144, 8),
     to_unsigned(145, 8),
     to_unsigned(146, 8),
     to_unsigned(147, 8),
     to_unsigned(148, 8),
     to_unsigned(149, 8),
     to_unsigned(150, 8),
     to_unsigned(151, 8),
     to_unsigned(152, 8),
     to_unsigned(153, 8),
     to_unsigned(154, 8),
     to_unsigned(155, 8),
     to_unsigned(156, 8),
     to_unsigned(157, 8),
     to_unsigned(158, 8),
     to_unsigned(159, 8));

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l288_c13_fe56_return_output;
     VAR_chacha20poly1305_decrypt_key := VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l183_l158_DUPLICATE_0a36_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_fbb8_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l150_c9_fbb8_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_cf38_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l149_c9_cf38_return_output;
     VAR_chacha20poly1305_decrypt_nonce := VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_f336_return_output;
     -- uint8_array32_be[chacha20poly1305_decrypt_tb_c_l183_c41_a342] LATENCY=0
     VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output := uint8_array32_be(
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l183_l158_DUPLICATE_0a36_return_output);

     -- uint8_array12_be[chacha20poly1305_decrypt_tb_c_l184_c40_1caa] LATENCY=0
     VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_1caa_return_output := uint8_array12_be(
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l159_l184_DUPLICATE_f336_return_output);

     -- Submodule level 2
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_1caa_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_1caa_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l184_c40_1caa_return_output;
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l183_c41_a342_return_output;
     -- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l183_c179_093b] LATENCY=0
     -- Inputs
     CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_x <= VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_x;
     -- Outputs
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output := CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l183_c302_1489] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output;

     -- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l183_c210_a1cc] LATENCY=0
     -- Inputs
     CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_x <= VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_x;
     -- Outputs
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output := CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l184_c130_4c71] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l183_c332_d4d8] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l184_c100_1c53] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output;

     -- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l183_c117_2a9b] LATENCY=0
     -- Inputs
     CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_x <= VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_x;
     -- Outputs
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output := CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output;

     -- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l183_c148_c11e] LATENCY=0
     -- Inputs
     CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_x <= VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_x;
     -- Outputs
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output := CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l183_c272_c1b2] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l184_c160_32aa] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l183_c241_1fac] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg0 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l184_c100_1c53_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg0 := resize(VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l183_c117_2a9b_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg4 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l183_c241_1fac_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg2 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l184_c160_32aa_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg7 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l183_c332_d4d8_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg3 := resize(VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l183_c210_a1cc_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg1 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l184_c130_4c71_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg1 := resize(VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l183_c148_c11e_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg5 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l183_c272_c1b2_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg2 := resize(VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l183_c179_093b_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg6 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l183_c302_1489_return_output, 32);
 -- Reads from global variables
     VAR_chacha20poly1305_decrypt_axis_in_ready := global_to_module.chacha20poly1305_decrypt_axis_in_ready;
     VAR_chacha20poly1305_decrypt_axis_out := global_to_module.chacha20poly1305_decrypt_axis_out;
     -- Submodule level 0
     VAR_return_output := VAR_chacha20poly1305_decrypt_axis_out;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_right := VAR_chacha20poly1305_decrypt_axis_in_ready;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg1 := resize(VAR_chacha20poly1305_decrypt_axis_in_ready, 32);
     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_3f2c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_3f2c_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(8);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_b684 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_b684_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(3);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_0801 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_0801_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(6);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_c83e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_c83e_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(0);

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d[chacha20poly1305_decrypt_tb_c_l251_c58_9d96] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l251_c58_9d96_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_36c1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_36c1_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(2);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d[chacha20poly1305_decrypt_tb_c_l248_c8_c79e] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l248_c8_c79e_return_output := VAR_chacha20poly1305_decrypt_axis_out.valid;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_7af8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_7af8_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(15);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_5abe LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_5abe_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(5);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_be47 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_be47_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(10);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_eac9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_eac9_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(7);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_a48c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_a48c_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(9);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_eeb6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_eeb6_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(13);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d[chacha20poly1305_decrypt_tb_c_l268_c12_928d] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tlast;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_37db LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_37db_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(1);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_ef83 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_ef83_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(11);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_671b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_671b_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(12);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_efbd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_efbd_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(4);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_8e59 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_8e59_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(14);

     -- Submodule level 1
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_efbd_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_efbd_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_c83e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_c83e_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_3f2c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_3f2c_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_7af8_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_7af8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_b684_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_b684_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_8e59_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_8e59_return_output, 32);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l268_c12_928d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_671b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_671b_return_output, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_left := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l248_c8_c79e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_a48c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_a48c_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_eac9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_eac9_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_ef83_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_ef83_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_be47_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_be47_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_eeb6_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_eeb6_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_37db_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_37db_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_0801_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_0801_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_36c1_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_DUPLICATE_36c1_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_5abe_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l258_l262_DUPLICATE_5abe_return_output;
     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l251_c41_5695] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l251_c41_5695_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l251_c58_9d96_return_output);

     -- Submodule level 2
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l251_c41_5695_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l251_c41_5695_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l251_c41_5695_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l251_c41_5695_return_output;
     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l251_c200_2176] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l251_c230_8416] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l251_c169_6c9e] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l251_c260_51b2] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l251_c230_8416_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l251_c169_6c9e_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l251_c260_51b2_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l251_c200_2176_return_output, 32);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iftrue := VAR_CLOCK_ENABLE;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse := ciphertext_in_stream;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse := ciphertext_remaining_in;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_left := cycle_counter;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_left := cycle_counter;
     VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_left := cycle_counter;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg0 := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_left := input_packet_count;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_var_dim_0 := resize(input_packet_count, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_var_dim_0 := resize(input_packet_count, 1);
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg0 := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_arg0 := input_packet_count;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_left := output_packet_count;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_left := output_packet_count;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_var_dim_0 := resize(output_packet_count, 1);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_var_dim_0 := resize(output_packet_count, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_arg0 := output_packet_count;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse := plaintext_out_expected;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse := plaintext_out_size;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse := plaintext_remaining_out;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse := tag_match_checked;
     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l248_c8_f415] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l194_c30_26c6] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l230_c12_c373] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l237_c17_bf36] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output;

     -- chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee(
     chacha20poly1305_decrypt_axis_in,
     to_unsigned(0, 1));

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l190_c35_6769] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output;

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l205_c9_1d2f] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l179_c8_09da] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l189_c32_0b54] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output;

     -- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l198_c34_97d4] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_0;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_ref_toks_1;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output := VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output;

     -- BIN_OP_MOD[chacha20poly1305_decrypt_tb_c_l205_c31_26fa] LATENCY=0
     -- Inputs
     BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_left <= VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_left;
     BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_right <= VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_right;
     -- Outputs
     VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output := BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l286_c41_a2b3] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l296_c9_e3e9] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l324_c5_e824] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l230_c12_c373_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l248_c8_f415_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l179_c8_09da_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_left := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c9_1d2f_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_right := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l286_c41_a2b3_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_left := VAR_BIN_OP_MOD_chacha20poly1305_decrypt_tb_c_l205_c31_26fa_return_output;
     VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l237_c17_6bb4 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l237_c17_bf36_return_output, 32);
     VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l296_c9_e3e9_return_output, 32);
     VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l324_c5_b8b3 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l324_c5_e824_return_output, 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c35_6769_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l194_c30_26c6_return_output;
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l198_c9_532c := VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c34_97d4_return_output.data;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l189_c9_b205 := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l189_c32_0b54_return_output.data;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l189_c9_b205;
     REG_VAR_cycle_counter := VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l324_c5_b8b3;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l237_c17_6bb4;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_right := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_left := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55, 1);
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg0 := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l296_c9_cf55;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l198_c9_532c;
     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l180_c1_7711] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l297_c12_2242] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;

     -- VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l311_c42_328d] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_0;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_ref_toks_1;
     VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output := VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l307_c38_317b] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l249_c1_f913] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l179_c5_2e6b] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l205_c31_15f7] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output;

     -- Submodule level 2
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_right := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l205_c31_15f7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l297_c12_2242_return_output;
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l180_c1_7711_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l249_c1_f913_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l307_c38_317b_return_output;
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l311_c17_860d := VAR_VAR_REF_RD_uint8_t_128_uint8_t_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l311_c42_328d_return_output.data;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_left := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_right := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output, 33)));
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_expr := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l311_c17_860d;
     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(143);

     -- CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(41);

     -- CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(62);

     -- CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(122);

     -- CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(20);

     -- CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(67);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(130);

     -- CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(11);

     -- CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(100);

     -- CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(73);

     -- CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(49);

     -- CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(126);

     -- CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(66);

     -- CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(63);

     -- CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(8);

     -- CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(20);

     -- UNARY_OP_NOT[chacha20poly1305_decrypt_tb_c_l286_c69_ef49] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_expr <= VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output := UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(108);

     -- CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(27);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(114);

     -- CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(53);

     -- CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(89);

     -- CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(38);

     -- CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(86);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(35);

     -- CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(56);

     -- CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(47);

     -- CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(101);

     -- CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(24);

     -- CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(60);

     -- CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(48);

     -- CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(24);

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l268_c1_2dea] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(55);

     -- CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(114);

     -- CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(102);

     -- CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(29);

     -- CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(37);

     -- CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(72);

     -- CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(41);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(103);

     -- CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(65);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(10);

     -- CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(97);

     -- CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(50);

     -- CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(36);

     -- CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(34);

     -- CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(127);

     -- CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(117);

     -- CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(61);

     -- CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(86);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(141);

     -- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l227_c56_6fd6] LATENCY=0
     -- Inputs
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_left <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_left;
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_right <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_right;
     -- Outputs
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output := BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(96);

     -- CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(69);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b[chacha20poly1305_decrypt_tb_c_l251_c105_b34b] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_chacha20poly1305_decrypt_tb_c_l251_c105_b34b_arg3;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(80);

     -- CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(84);

     -- CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(28);

     -- print_aad[chacha20poly1305_decrypt_tb_c_l185_c9_3334] LATENCY=0
     -- Clock enable
     print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_CLOCK_ENABLE <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_CLOCK_ENABLE;
     -- Inputs
     print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad;
     print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad_len <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l185_c9_3334_aad_len;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(64);

     -- CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(52);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(140);

     -- CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(81);

     -- CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(103);

     -- CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(7);

     -- CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(59);

     -- CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(75);

     -- CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(74);

     -- CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(27);

     -- CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(30);

     -- CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(108);

     -- CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(105);

     -- CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(3);

     -- CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(93);

     -- CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(25);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(126);

     -- CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(39);

     -- CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(99);

     -- CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(111);

     -- CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(80);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(117);

     -- CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(58);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(135);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(120);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(128);

     -- CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(54);

     -- CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(110);

     -- CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(102);

     -- CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(109);

     -- CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(85);

     -- CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(98);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(119);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(127);

     -- CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(79);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(115);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(112);

     -- CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(22);

     -- CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(77);

     -- CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(4);

     -- CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(45);

     -- CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(76);

     -- CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(101);

     -- CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(16);

     -- CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(68);

     -- CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(92);

     -- printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165[chacha20poly1305_decrypt_tb_c_l181_c9_9165] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l181_c9_9165_chacha20poly1305_decrypt_tb_c_l181_c9_9165_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(72);

     -- CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(95);

     -- CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(12);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(68);

     -- CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(79);

     -- CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(61);

     -- CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(95);

     -- CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(97);

     -- CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(82);

     -- CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(32);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(138);

     -- CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(76);

     -- CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(83);

     -- CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(93);

     -- CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(67);

     -- CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(10);

     -- CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(46);

     -- CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(19);

     -- CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(70);

     -- CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(100);

     -- CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(23);

     -- CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(16);

     -- CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(31);

     -- CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(58);

     -- CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(104);

     -- CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(57);

     -- CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(94);

     -- CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(29);

     -- CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(83);

     -- CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(36);

     -- CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(75);

     -- CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(14);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l279_c17_fb4e] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(15);

     -- CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(96);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(137);

     -- CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(85);

     -- CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(55);

     -- CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(84);

     -- CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(59);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(118);

     -- CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(71);

     -- CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(90);

     -- CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(5);

     -- CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(35);

     -- CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(123);

     -- CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(6);

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l276_c16_9117] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(104);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(132);

     -- CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(52);

     -- CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(78);

     -- CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(7);

     -- CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(53);

     -- CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(106);

     -- CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(66);

     -- CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(40);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(1);

     -- CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(2);

     -- CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(18);

     -- CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(43);

     -- CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(3);

     -- CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(43);

     -- CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(21);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(39);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(105);

     -- CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(17);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(116);

     -- CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(74);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(120);

     -- CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(64);

     -- CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(13);

     -- CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(91);

     -- CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(88);

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l275_c1_88c6] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(107);

     -- CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(4);

     -- CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(94);

     -- CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(44);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(131);

     -- CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(63);

     -- CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(50);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(129);

     -- CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(121);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(25);

     -- CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(49);

     -- CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(98);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(113);

     -- CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(88);

     -- CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(115);

     -- CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(11);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(0);

     -- CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(26);

     -- CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(18);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(119);

     -- CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(33);

     -- CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(21);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(122);

     -- CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(26);

     -- CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(28);

     -- CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(69);

     -- CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(23);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(99);

     -- CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(30);

     -- CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(92);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l269_c16_4da1] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(125);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(142);

     -- CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(9);

     -- CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(57);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(124);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(139);

     -- CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(56);

     -- CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(116);

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l205_c9_cfd1] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(54);

     -- CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(82);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(62);

     -- CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(5);

     -- CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(37);

     -- CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(1);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(134);

     -- CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(77);

     -- CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(107);

     -- CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(110);

     -- CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(44);

     -- CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(73);

     -- CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(106);

     -- CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(13);

     -- CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(32);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(91);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(136);

     -- CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(48);

     -- CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(87);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(60);

     -- CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(111);

     -- CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(6);

     -- printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1[chacha20poly1305_decrypt_tb_c_l184_c65_d1b1] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_chacha20poly1305_decrypt_tb_c_l184_c65_d1b1_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(123);

     -- CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(22);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(78);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d[chacha20poly1305_decrypt_tb_c_l240_c173_7af9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(133);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(113);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_left <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_left;
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_right <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output := BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(51);

     -- CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(40);

     -- CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(118);

     -- printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743[chacha20poly1305_decrypt_tb_c_l183_c64_5743] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg3;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg4 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg4;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg5 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg5;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg6 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg6;
     printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg7 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l183_c64_5743_chacha20poly1305_decrypt_tb_c_l183_c64_5743_arg7;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(14);

     -- CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(42);

     -- CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(71);

     -- CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(65);

     -- CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(42);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(121);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l213_c8_7e08] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(38);

     -- FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d[chacha20poly1305_decrypt_tb_c_l280_c168_de5e] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(125);

     -- CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(8);

     -- CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(45);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(33);

     -- CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(109);

     -- CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(70);

     -- printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0[chacha20poly1305_decrypt_tb_c_l191_c9_8ae0] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_chacha20poly1305_decrypt_tb_c_l191_c9_8ae0_arg1;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(0);

     -- CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(51);

     -- CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(112);

     -- CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(31);

     -- CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(17);

     -- CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(90);

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l221_c16_e55e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_left;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(87);

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l256_c16_8247] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(9);

     -- CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(46);

     -- CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(89);

     -- CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(19);

     -- CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(12);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l239_c17_0476] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(34);

     -- CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(15);

     -- CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(2);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l205_c59_fd85] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(47);

     -- CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(124);

     -- printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0[chacha20poly1305_decrypt_tb_c_l200_c9_53d0] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_chacha20poly1305_decrypt_tb_c_l200_c9_53d0_arg1;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output(81);

     -- Submodule level 3
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_left := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_cfd1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l276_c16_9117_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_right := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l205_c59_fd85_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l213_c8_7e08_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l269_c16_4da1_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l239_c17_0476_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l279_c17_fb4e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l260_DUPLICATE_714c_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output, 32);
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_0_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_66f7_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_100_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_031d_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_101_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_decf_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_102_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_4c3e_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_103_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_16d9_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_104_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_81a1_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_105_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_7cdc_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_106_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_d349_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_107_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_108_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_8329_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_109_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_1e0f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output, 32);
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_10_d41d_chacha20poly1305_decrypt_tb_c_l262_l258_l276_l248_l268_DUPLICATE_932c_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_110_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_b9bf_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_111_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3394_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output, 32);
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l276_l258_DUPLICATE_8759_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output, 32);
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_12_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_70ac_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output, 32);
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l262_l258_l276_DUPLICATE_1fa2_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output, 32);
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_14_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l262_l248_l268_DUPLICATE_f117_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output, 32);
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_15_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_a798_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_16_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5e58_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_17_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_4744_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_18_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6c59_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_19_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_7555_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output, 32);
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_1_d41d_chacha20poly1305_decrypt_tb_c_l276_l262_l248_l268_l258_DUPLICATE_17f7_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_20_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_940d_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_21_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_b4c4_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_22_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_e56c_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_23_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_71a2_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_24_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_3653_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_25_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_f12b_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_26_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_73cd_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_27_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_38bc_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_28_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_43b9_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_29_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_1855_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output, 32);
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_2_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_7070_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_30_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_3850_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_31_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_ff54_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_32_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5403_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_33_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_ff42_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_34_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_f654_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_35_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l248_l276_DUPLICATE_78f5_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_36_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_9dc4_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_37_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_1d2d_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_38_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_fe6f_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_39_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_d22e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output, 32);
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l268_l258_l276_DUPLICATE_d0cc_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_40_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_9192_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_41_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_2c70_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_42_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_317f_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_43_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_628b_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_44_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_2c59_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_45_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a9bc_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_46_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l248_l276_DUPLICATE_f267_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_47_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_0e0a_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_48_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_be6e_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_49_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_ecd4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output, 32);
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_4_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_fe15_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_50_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_d365_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_51_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_f1ef_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_52_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4e13_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_53_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l268_l248_DUPLICATE_5bab_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_54_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_fe01_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_55_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_1b2c_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_56_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_1eba_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_57_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_2864_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_58_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_114a_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_59_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l268_l276_DUPLICATE_a634_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output, 32);
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_5_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l268_l258_l276_DUPLICATE_5cf2_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_60_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_6561_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_61_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l280_l248_DUPLICATE_48e0_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_62_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l276_l280_DUPLICATE_b262_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_63_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_09c9_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_64_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_040f_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_65_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_7743_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_66_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_4c60_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_67_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_e6c0_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_68_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_1e52_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_69_d41d_chacha20poly1305_decrypt_tb_c_l276_l280_l248_l268_DUPLICATE_bd12_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output, 32);
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_6_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l268_l258_l248_DUPLICATE_9dca_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_70_d41d_chacha20poly1305_decrypt_tb_c_l276_l268_l248_l280_DUPLICATE_91d8_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_71_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l280_l276_DUPLICATE_5c1a_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_72_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_3506_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_73_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_e356_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_74_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_a199_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_75_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_cfe7_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_76_d41d_chacha20poly1305_decrypt_tb_c_l248_l268_l280_l276_DUPLICATE_be83_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_77_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_7c0f_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_78_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_1ebf_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_79_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l276_l268_DUPLICATE_50bb_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output, 32);
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_7_d41d_chacha20poly1305_decrypt_tb_c_l276_l258_l248_l268_l262_DUPLICATE_128f_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_80_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_97d8_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_81_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l268_l280_DUPLICATE_9da9_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_82_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_6566_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_83_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_528d_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_84_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_0852_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_85_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_0727_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_86_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_9a7d_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_87_d41d_chacha20poly1305_decrypt_tb_c_l268_l248_l276_l280_DUPLICATE_f275_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_88_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_9425_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_89_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l248_l280_DUPLICATE_63da_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output, 32);
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_8_d41d_chacha20poly1305_decrypt_tb_c_l262_l276_l258_l248_l268_DUPLICATE_e896_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_90_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_c6ae_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_91_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_2513_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_92_d41d_chacha20poly1305_decrypt_tb_c_l248_l276_l268_l280_DUPLICATE_abe2_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_93_d41d_chacha20poly1305_decrypt_tb_c_l248_l280_l268_l276_DUPLICATE_5c64_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_94_d41d_chacha20poly1305_decrypt_tb_c_l276_l248_l280_l268_DUPLICATE_5468_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_95_d41d_chacha20poly1305_decrypt_tb_c_l280_l248_l276_l268_DUPLICATE_e9be_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_96_d41d_chacha20poly1305_decrypt_tb_c_l280_l268_l276_l248_DUPLICATE_e11b_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_97_d41d_chacha20poly1305_decrypt_tb_c_l268_l276_l280_l248_DUPLICATE_cc73_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_98_d41d_chacha20poly1305_decrypt_tb_c_l268_l280_l276_l248_DUPLICATE_6c92_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_99_d41d_chacha20poly1305_decrypt_tb_c_l280_l276_l248_l268_DUPLICATE_baf5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 := resize(VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output, 32);
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_128_9_d41d_chacha20poly1305_decrypt_tb_c_l258_l276_l248_l262_l268_DUPLICATE_ff7a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_53e7_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_c86e_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_04b9_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_834f_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_9e7c_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_8696_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_5029_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_dfbc_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_15d7_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5610_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_7cbf_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l223_l234_l213_l230_DUPLICATE_5ff1_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_738e_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_6844_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2de5_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l240_l230_DUPLICATE_da77_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_162c_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_afc4_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_fdcf_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_b2eb_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_edfa_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_75a7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l223_DUPLICATE_a439_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_cbdf_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_7e23_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_3df8_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_6c82_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1f7d_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_124b_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_d35b_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l240_l234_DUPLICATE_e9d7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_3537_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l223_DUPLICATE_3b63_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_6e02_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l213_l230_DUPLICATE_0464_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_e478_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_e817_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_24a0_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_1e64_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_c7b3_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_5295_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_f618_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_66e1_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_2b6f_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_fa4b_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_92a8_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_c75f_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_f3d8_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_788a_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_556b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l223_l213_l234_l230_DUPLICATE_e16c_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_ea10_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_4e76_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_918e_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_f518_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l230_l240_DUPLICATE_9e4b_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_85c7_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_8bd7_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_b4c9_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_966b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_fe75_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_167a_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_e855_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_9978_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_90f1_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_642c_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_2020_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_1588_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_2c1d_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_280c_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l240_DUPLICATE_9249_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l223_DUPLICATE_6e39_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_dc64_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_cdb3_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_5890_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_9704_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l213_l230_l234_l240_DUPLICATE_9bc2_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_028d_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_4ed8_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_16a2_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_82a4_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_bfcf_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l213_l223_DUPLICATE_29b3_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2dbf_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_67e0_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l234_l240_l230_l213_DUPLICATE_e7b0_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_82ac_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_e537_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_b293_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_0661_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l234_l230_DUPLICATE_d097_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_5f5d_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l230_l213_DUPLICATE_b384_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l223_l234_DUPLICATE_313b_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_5e01_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_591e_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l234_l213_DUPLICATE_e646_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_72f3_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_c6e8_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_dfd5_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_bb66_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_ca42_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_fd37_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l230_l234_DUPLICATE_1edc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l230_l223_l213_l234_DUPLICATE_323c_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_89a0_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_8f64_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_572c_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l230_l234_l240_l213_DUPLICATE_0289_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l234_l213_l230_l240_DUPLICATE_686f_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_72ad_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l240_l234_DUPLICATE_d660_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_bb93_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_bcda_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_1ed4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l234_l223_l230_l213_DUPLICATE_183c_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l240_l234_l213_l230_DUPLICATE_a386_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l240_l213_DUPLICATE_7b2c_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l213_l240_l230_l234_DUPLICATE_3671_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_1811_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l230_l240_l213_l234_DUPLICATE_be20_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l240_l213_l234_l230_DUPLICATE_b2c2_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l213_l234_l240_l230_DUPLICATE_ec0c_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l234_l230_l213_l240_DUPLICATE_99cf_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l240_l230_l213_l234_DUPLICATE_f526_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l230_l213_l234_l240_DUPLICATE_2e2d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l223_l230_l213_l234_DUPLICATE_97cd_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_88c6_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l221_c16_e55e_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c46_2515_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l240_c173_7af9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l256_c16_8247_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_100_CONST_REF_RD_uint8_t_uint8_t_128_116_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_101_CONST_REF_RD_uint8_t_uint8_t_128_117_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_102_CONST_REF_RD_uint8_t_uint8_t_128_118_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_103_CONST_REF_RD_uint8_t_uint8_t_128_119_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_104_CONST_REF_RD_uint8_t_uint8_t_128_120_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_105_CONST_REF_RD_uint8_t_uint8_t_128_121_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_106_CONST_REF_RD_uint8_t_uint8_t_128_122_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_107_CONST_REF_RD_uint8_t_uint8_t_128_123_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_108_CONST_REF_RD_uint8_t_uint8_t_128_124_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_109_CONST_REF_RD_uint8_t_uint8_t_128_125_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_110_CONST_REF_RD_uint8_t_uint8_t_128_126_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_111_CONST_REF_RD_uint8_t_uint8_t_128_127_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_96_CONST_REF_RD_uint8_t_uint8_t_128_112_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_97_CONST_REF_RD_uint8_t_uint8_t_128_113_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_98_CONST_REF_RD_uint8_t_uint8_t_128_114_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l280_c46_919e_ITER_99_CONST_REF_RD_uint8_t_uint8_t_128_115_d41d_chacha20poly1305_decrypt_tb_c_l280_c168_de5e_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l268_c1_2dea_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_right := VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l286_c69_ef49_return_output;
     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l214_c1_8bf9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l269_c13_ea14] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l269_c1_5c29] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l205_c9_2fad] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l271_c1_bc29] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l276_c1_6034] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_d75f] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l221_c13_8dac] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output := FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l234_c13_8907] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l260_c47_e8d9] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l276_c13_7c6a] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l258_c20_b069] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_left;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;

     -- Submodule level 4
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l205_c9_2fad_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l271_c1_bc29_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l258_c20_b069_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l260_c47_e8d9_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_d75f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l214_c1_8bf9_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l269_c1_5c29_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l276_c1_6034_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l234_c13_8907_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l269_c13_ea14_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l276_c13_7c6a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l260_c30_1002_0;
     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed[chacha20poly1305_decrypt_tb_c_l232_c62_514c] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l232_c62_514c_return_output := CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed(
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output);

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l231_c1_de39] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d[chacha20poly1305_decrypt_tb_c_l277_c18_784d] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l277_c18_784d_chacha20poly1305_decrypt_tb_c_l277_c18_784d_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l205_c1_c273] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b[chacha20poly1305_decrypt_tb_c_l272_c17_fb9b] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_chacha20poly1305_decrypt_tb_c_l272_c17_fb9b_arg0;
     -- Outputs

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c(
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l217_c9_f138_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l221_c13_8dac_return_output,
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l227_c56_6fd6_return_output,
     to_unsigned(1, 1));

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l259_c1_58ca] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output := FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd[chacha20poly1305_decrypt_tb_c_l270_c17_aafd] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_chacha20poly1305_decrypt_tb_c_l270_c17_aafd_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l230_c9_1787] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l268_c9_cfd7] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;

     -- Submodule level 5
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l259_c1_58ca_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l205_c1_c273_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l231_c1_de39_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l230_c9_1787_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l268_c9_cfd7_return_output;
     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l234_c1_b6b6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68[chacha20poly1305_decrypt_tb_c_l206_c9_6d68] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_chacha20poly1305_decrypt_tb_c_l206_c9_6d68_arg1;
     -- Outputs

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l232_c45_3245] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l232_c45_3245_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l232_c62_514c_return_output);

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f[chacha20poly1305_decrypt_tb_c_l261_c21_a17f] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l254_c9_d8d6_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_chacha20poly1305_decrypt_tb_c_l261_c21_a17f_arg2;
     -- Outputs

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l213_c5_1de4] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l248_c5_da03] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;

     -- Submodule level 6
     VAR_printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l234_c1_b6b6_return_output;
     REG_VAR_chacha20poly1305_decrypt_axis_in := VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_left := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_left := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_var_dim_0 := resize(VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_var_dim_0 := resize(VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output, 1);
     REG_VAR_input_packet_count := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg0 := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l232_c45_3245_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l232_c45_3245_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l232_c45_3245_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l232_c45_3245_return_output;
     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l232_c267_3cbf] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d[chacha20poly1305_decrypt_tb_c_l235_c17_7f1d] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_chacha20poly1305_decrypt_tb_c_l235_c17_7f1d_arg0;
     -- Outputs

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l232_c207_f310] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output;

     -- CONST_REF_RD_uint8_t_128_uint8_t_128_7166_chacha20poly1305_decrypt_tb_c_l297_l286_l300_DUPLICATE_f22f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_7166_chacha20poly1305_decrypt_tb_c_l297_l286_l300_DUPLICATE_f22f_return_output := CONST_REF_RD_uint8_t_128_uint8_t_128_7166(
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output,
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l248_c5_da03_return_output);

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l232_c176_e3c5] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l300_c17_b9d8] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l302_c40_0822] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output;

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6_chacha20poly1305_decrypt_tb_c_l286_l300_l297_DUPLICATE_55b0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6_chacha20poly1305_decrypt_tb_c_l286_l300_l297_DUPLICATE_55b0_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6(
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l179_c5_2e6b_return_output,
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output,
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l213_c5_1de4_return_output);

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l232_c237_0c4e] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l286_c9_4b3b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l303_c43_94e2] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output;

     -- Submodule level 7
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_left := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c9_4b3b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l300_c17_b9d8_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_7166_chacha20poly1305_decrypt_tb_c_l297_l286_l300_DUPLICATE_f22f_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse := VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_7166_chacha20poly1305_decrypt_tb_c_l297_l286_l300_DUPLICATE_f22f_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse := VAR_CONST_REF_RD_uint8_t_128_uint8_t_128_7166_chacha20poly1305_decrypt_tb_c_l297_l286_l300_DUPLICATE_f22f_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6_chacha20poly1305_decrypt_tb_c_l286_l300_l297_DUPLICATE_55b0_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6_chacha20poly1305_decrypt_tb_c_l286_l300_l297_DUPLICATE_55b0_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_d1f6_chacha20poly1305_decrypt_tb_c_l286_l300_l297_DUPLICATE_55b0_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l232_c267_3cbf_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l232_c237_0c4e_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l232_c207_f310_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l232_c176_e3c5_return_output, 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l303_c43_94e2_return_output;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l302_c17_010b := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l302_c40_0822_return_output.data;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l302_c17_010b;
     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l286_c9_e09e] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l300_c13_23ed] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1[chacha20poly1305_decrypt_tb_c_l232_c108_5fc1] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_chacha20poly1305_decrypt_tb_c_l232_c108_5fc1_arg3;
     -- Outputs

     -- Submodule level 8
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_left := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_e09e_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l300_c13_23ed_return_output;
     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l286_c9_21ab] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l297_c9_b19f] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;

     -- Submodule level 9
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l286_c9_21ab_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l297_c9_b19f_return_output;
     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l287_c1_acb3] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l286_c5_dbd1] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;

     -- Submodule level 10
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l287_c1_acb3_return_output;
     REG_VAR_ciphertext_in_stream := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     REG_VAR_ciphertext_remaining_in := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_right := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     REG_VAR_output_packet_count := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     REG_VAR_plaintext_out_expected := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     REG_VAR_plaintext_out_size := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     REG_VAR_plaintext_remaining_out := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iffalse := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l286_c5_dbd1_return_output;
     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l291_c1_cbc7] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l289_c1_ec75] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output;

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l320_c9_eb04] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l298_c1_84a2] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output;

     -- Submodule level 11
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l320_c9_eb04_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l291_c1_cbc7_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l289_c1_ec75_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l298_c1_84a2_return_output;
     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l320_c5_c1e4] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l300_c1_bafe] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695[chacha20poly1305_decrypt_tb_c_l290_c13_9695] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c13_9695_chacha20poly1305_decrypt_tb_c_l290_c13_9695_arg0;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a[chacha20poly1305_decrypt_tb_c_l292_c13_395a] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l292_c13_395a_chacha20poly1305_decrypt_tb_c_l292_c13_395a_arg0;
     -- Outputs

     -- Submodule level 12
     VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l300_c1_bafe_return_output;
     REG_VAR_tag_match_checked := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l320_c5_c1e4_return_output;
     -- printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4[chacha20poly1305_decrypt_tb_c_l304_c17_01e4] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_chacha20poly1305_decrypt_tb_c_l304_c17_01e4_arg1;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e[chacha20poly1305_decrypt_tb_c_l313_c17_391e] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l313_c17_391e_chacha20poly1305_decrypt_tb_c_l313_c17_391e_arg1;
     -- Outputs

     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_input_packet_count <= REG_VAR_input_packet_count;
REG_COMB_ciphertext_in_stream <= REG_VAR_ciphertext_in_stream;
REG_COMB_ciphertext_remaining_in <= REG_VAR_ciphertext_remaining_in;
REG_COMB_cycle_counter <= REG_VAR_cycle_counter;
REG_COMB_output_packet_count <= REG_VAR_output_packet_count;
REG_COMB_plaintext_out_size <= REG_VAR_plaintext_out_size;
REG_COMB_plaintext_remaining_out <= REG_VAR_plaintext_remaining_out;
REG_COMB_plaintext_out_expected <= REG_VAR_plaintext_out_expected;
REG_COMB_tag_match_checked <= REG_VAR_tag_match_checked;
REG_COMB_chacha20poly1305_decrypt_axis_in <= REG_VAR_chacha20poly1305_decrypt_axis_in;
-- Global wires driven various places in pipeline
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_key <= VAR_chacha20poly1305_decrypt_key;
else
  module_to_global.chacha20poly1305_decrypt_key <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_nonce <= VAR_chacha20poly1305_decrypt_nonce;
else
  module_to_global.chacha20poly1305_decrypt_nonce <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad <= VAR_chacha20poly1305_decrypt_aad;
else
  module_to_global.chacha20poly1305_decrypt_aad <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad_len <= VAR_chacha20poly1305_decrypt_aad_len;
else
  module_to_global.chacha20poly1305_decrypt_aad_len <= to_unsigned(0, 8);
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= VAR_chacha20poly1305_decrypt_axis_out_ready;
else
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= to_unsigned(0, 1);
end if;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     input_packet_count <= REG_COMB_input_packet_count;
     ciphertext_in_stream <= REG_COMB_ciphertext_in_stream;
     ciphertext_remaining_in <= REG_COMB_ciphertext_remaining_in;
     cycle_counter <= REG_COMB_cycle_counter;
     output_packet_count <= REG_COMB_output_packet_count;
     plaintext_out_size <= REG_COMB_plaintext_out_size;
     plaintext_remaining_out <= REG_COMB_plaintext_remaining_out;
     plaintext_out_expected <= REG_COMB_plaintext_out_expected;
     tag_match_checked <= REG_COMB_tag_match_checked;
     chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in;
 end if;
 end if;
end process;
-- Shared global regs
module_to_global.chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in when clk_en_internal='1' else chacha20poly1305_decrypt_axis_in;

end arch;
