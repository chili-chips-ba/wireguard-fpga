mem['h0000] = 32'h00001517;
mem['h0001] = 32'h08C50513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'h00860613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFE850513;
mem['h000E] = 32'h10001597;
mem['h000F] = 32'h3F458593;
mem['h0010] = 32'h00B55863;
mem['h0011] = 32'h00052023;
mem['h0012] = 32'h00450513;
mem['h0013] = 32'hFEB54CE3;
mem['h0014] = 32'h10008117;
mem['h0015] = 32'hFB010113;
mem['h0016] = 32'h10000197;
mem['h0017] = 32'h7C018193;
mem['h0018] = 32'h00A54533;
mem['h0019] = 32'h00B5C5B3;
mem['h001A] = 32'h00C64633;
mem['h001B] = 32'h48C000EF;
mem['h001C] = 32'h0000006F;
mem['h001D] = 32'h00452783;
mem['h001E] = 32'h0087A783;
mem['h001F] = 32'h0007A783;
mem['h0020] = 32'h0007A783;
mem['h0021] = 32'hFE07C8E3;
mem['h0022] = 32'h00452783;
mem['h0023] = 32'h0087A783;
mem['h0024] = 32'h0007A783;
mem['h0025] = 32'h00B78023;
mem['h0026] = 32'h00008067;
mem['h0027] = 32'hFE010113;
mem['h0028] = 32'h00812C23;
mem['h0029] = 32'h01212823;
mem['h002A] = 32'hFFF60413;
mem['h002B] = 32'h00001937;
mem['h002C] = 32'h00912A23;
mem['h002D] = 32'h01312623;
mem['h002E] = 32'h00112E23;
mem['h002F] = 32'h00050493;
mem['h0030] = 32'h00058993;
mem['h0031] = 32'h00241413;
mem['h0032] = 32'hEE890913;
mem['h0033] = 32'h0089D7B3;
mem['h0034] = 32'h00F7F793;
mem['h0035] = 32'h00F907B3;
mem['h0036] = 32'h0007C583;
mem['h0037] = 32'h00048513;
mem['h0038] = 32'hFFC40413;
mem['h0039] = 32'hF91FF0EF;
mem['h003A] = 32'hFE0452E3;
mem['h003B] = 32'h01C12083;
mem['h003C] = 32'h01812403;
mem['h003D] = 32'h01412483;
mem['h003E] = 32'h01012903;
mem['h003F] = 32'h00C12983;
mem['h0040] = 32'h02010113;
mem['h0041] = 32'h00008067;
mem['h0042] = 32'h0A058863;
mem['h0043] = 32'hFE010113;
mem['h0044] = 32'h00912A23;
mem['h0045] = 32'h00058493;
mem['h0046] = 32'h01312623;
mem['h0047] = 32'h00A00593;
mem['h0048] = 32'h00050993;
mem['h0049] = 32'h00048513;
mem['h004A] = 32'h00812C23;
mem['h004B] = 32'h00112E23;
mem['h004C] = 32'h01212823;
mem['h004D] = 32'h01412423;
mem['h004E] = 32'h505000EF;
mem['h004F] = 32'h0FF57513;
mem['h0050] = 32'h00100413;
mem['h0051] = 32'h06857E63;
mem['h0052] = 32'h00900A13;
mem['h0053] = 32'h00040593;
mem['h0054] = 32'h00048513;
mem['h0055] = 32'h4E9000EF;
mem['h0056] = 32'h0FF57913;
mem['h0057] = 32'h03090593;
mem['h0058] = 32'h0FF5F593;
mem['h0059] = 32'h00098513;
mem['h005A] = 32'hF0DFF0EF;
mem['h005B] = 32'h00040593;
mem['h005C] = 32'h00090513;
mem['h005D] = 32'h49D000EF;
mem['h005E] = 32'h40A487B3;
mem['h005F] = 32'h00A00593;
mem['h0060] = 32'h00040513;
mem['h0061] = 32'h0FF7F493;
mem['h0062] = 32'h00040913;
mem['h0063] = 32'h4B1000EF;
mem['h0064] = 32'h00050413;
mem['h0065] = 32'hFB2A6CE3;
mem['h0066] = 32'h01C12083;
mem['h0067] = 32'h01812403;
mem['h0068] = 32'h01412483;
mem['h0069] = 32'h01012903;
mem['h006A] = 32'h00C12983;
mem['h006B] = 32'h00812A03;
mem['h006C] = 32'h02010113;
mem['h006D] = 32'h00008067;
mem['h006E] = 32'h03000593;
mem['h006F] = 32'hEB9FF06F;
mem['h0070] = 32'h00241793;
mem['h0071] = 32'h00878433;
mem['h0072] = 32'h00141413;
mem['h0073] = 32'hF79FF06F;
mem['h0074] = 32'hFF010113;
mem['h0075] = 32'h00812423;
mem['h0076] = 32'h00912223;
mem['h0077] = 32'h00112623;
mem['h0078] = 32'h00050493;
mem['h0079] = 32'h00058413;
mem['h007A] = 32'h00044583;
mem['h007B] = 32'h00059C63;
mem['h007C] = 32'h00C12083;
mem['h007D] = 32'h00812403;
mem['h007E] = 32'h00412483;
mem['h007F] = 32'h01010113;
mem['h0080] = 32'h00008067;
mem['h0081] = 32'h00048513;
mem['h0082] = 32'h00140413;
mem['h0083] = 32'hE69FF0EF;
mem['h0084] = 32'hFD9FF06F;
mem['h0085] = 32'hFF010113;
mem['h0086] = 32'h00112623;
mem['h0087] = 32'h00812423;
mem['h0088] = 32'h00912223;
mem['h0089] = 32'h00058493;
mem['h008A] = 32'h0005C583;
mem['h008B] = 32'h00050413;
mem['h008C] = 32'hED9FF0EF;
mem['h008D] = 32'h00040513;
mem['h008E] = 32'h02E00593;
mem['h008F] = 32'hE39FF0EF;
mem['h0090] = 32'h0014C583;
mem['h0091] = 32'h00040513;
mem['h0092] = 32'hEC1FF0EF;
mem['h0093] = 32'h00040513;
mem['h0094] = 32'h02E00593;
mem['h0095] = 32'hE21FF0EF;
mem['h0096] = 32'h0024C583;
mem['h0097] = 32'h00040513;
mem['h0098] = 32'hEA9FF0EF;
mem['h0099] = 32'h00040513;
mem['h009A] = 32'h02E00593;
mem['h009B] = 32'hE09FF0EF;
mem['h009C] = 32'h00040513;
mem['h009D] = 32'h00812403;
mem['h009E] = 32'h0034C583;
mem['h009F] = 32'h00C12083;
mem['h00A0] = 32'h00412483;
mem['h00A1] = 32'h01010113;
mem['h00A2] = 32'hE81FF06F;
mem['h00A3] = 32'h100016B7;
mem['h00A4] = 32'h4286A703;
mem['h00A5] = 32'h100017B7;
mem['h00A6] = 32'hC2878793;
mem['h00A7] = 32'h00F707B3;
mem['h00A8] = 32'h00A70733;
mem['h00A9] = 32'h42E6A423;
mem['h00AA] = 32'h000016B7;
mem['h00AB] = 32'h80068693;
mem['h00AC] = 32'h00E6D463;
mem['h00AD] = 32'h00100073;
mem['h00AE] = 32'h00078513;
mem['h00AF] = 32'h00008067;
mem['h00B0] = 32'h00000793;
mem['h00B1] = 32'h00F58733;
mem['h00B2] = 32'h00074683;
mem['h00B3] = 32'h00F50733;
mem['h00B4] = 32'h00178793;
mem['h00B5] = 32'h00D70023;
mem['h00B6] = 32'hFEC796E3;
mem['h00B7] = 32'h00008067;
mem['h00B8] = 32'h00052783;
mem['h00B9] = 32'h0007A783;
mem['h00BA] = 32'h0187A783;
mem['h00BB] = 32'h0007A783;
mem['h00BC] = 32'h0007A783;
mem['h00BD] = 32'h0017F793;
mem['h00BE] = 32'h1E078E63;
mem['h00BF] = 32'h00052783;
mem['h00C0] = 32'h0005C703;
mem['h00C1] = 32'hFFFF8637;
mem['h00C2] = 32'h0007A783;
mem['h00C3] = 32'h00777713;
mem['h00C4] = 32'hFFFF08B7;
mem['h00C5] = 32'h0107A783;
mem['h00C6] = 32'hFFF60613;
mem['h00C7] = 32'h0007A683;
mem['h00C8] = 32'h0006A783;
mem['h00C9] = 32'hFF87F793;
mem['h00CA] = 32'h00E7E7B3;
mem['h00CB] = 32'h00F6A023;
mem['h00CC] = 32'h00052783;
mem['h00CD] = 32'h0015C703;
mem['h00CE] = 32'h0007A783;
mem['h00CF] = 32'h00777713;
mem['h00D0] = 32'h00371713;
mem['h00D1] = 32'h0107A783;
mem['h00D2] = 32'h0007A683;
mem['h00D3] = 32'h0006A783;
mem['h00D4] = 32'hFC77F793;
mem['h00D5] = 32'h00E7E7B3;
mem['h00D6] = 32'h00F6A023;
mem['h00D7] = 32'h00052783;
mem['h00D8] = 32'h0025C703;
mem['h00D9] = 32'h0007A783;
mem['h00DA] = 32'h00177713;
mem['h00DB] = 32'h00671713;
mem['h00DC] = 32'h0107A783;
mem['h00DD] = 32'h0007A683;
mem['h00DE] = 32'h0006A783;
mem['h00DF] = 32'hFBF7F793;
mem['h00E0] = 32'h00E7E7B3;
mem['h00E1] = 32'h00F6A023;
mem['h00E2] = 32'h00052783;
mem['h00E3] = 32'h0035C703;
mem['h00E4] = 32'h0007A783;
mem['h00E5] = 32'h00177713;
mem['h00E6] = 32'h00771713;
mem['h00E7] = 32'h0107A783;
mem['h00E8] = 32'h0007A683;
mem['h00E9] = 32'h0006A783;
mem['h00EA] = 32'hF7F7F793;
mem['h00EB] = 32'h00E7E7B3;
mem['h00EC] = 32'h00F6A023;
mem['h00ED] = 32'h00858713;
mem['h00EE] = 32'h00000793;
mem['h00EF] = 32'h00052683;
mem['h00F0] = 32'h00072803;
mem['h00F1] = 32'h01078793;
mem['h00F2] = 32'h0006A683;
mem['h00F3] = 32'h01070713;
mem['h00F4] = 32'h0006A683;
mem['h00F5] = 32'h0006A683;
mem['h00F6] = 32'h0106A023;
mem['h00F7] = 32'h00052683;
mem['h00F8] = 32'hFF472803;
mem['h00F9] = 32'h0006A683;
mem['h00FA] = 32'h0046A683;
mem['h00FB] = 32'h0006A683;
mem['h00FC] = 32'h0106A023;
mem['h00FD] = 32'h00052683;
mem['h00FE] = 32'hFF872803;
mem['h00FF] = 32'h0006A683;
mem['h0100] = 32'h0086A683;
mem['h0101] = 32'h0006A683;
mem['h0102] = 32'h0106A023;
mem['h0103] = 32'h00052683;
mem['h0104] = 32'hFFC72803;
mem['h0105] = 32'h0006A683;
mem['h0106] = 32'h00C6A683;
mem['h0107] = 32'h0006A683;
mem['h0108] = 32'h0106A023;
mem['h0109] = 32'h0045A683;
mem['h010A] = 32'h04D7FE63;
mem['h010B] = 32'h00052683;
mem['h010C] = 32'h0006A683;
mem['h010D] = 32'h0106A683;
mem['h010E] = 32'h0006A803;
mem['h010F] = 32'h00082683;
mem['h0110] = 32'h0116E6B3;
mem['h0111] = 32'h00D82023;
mem['h0112] = 32'h00052683;
mem['h0113] = 32'h0006A683;
mem['h0114] = 32'h0106A683;
mem['h0115] = 32'h0006A803;
mem['h0116] = 32'h00082683;
mem['h0117] = 32'h00C6F6B3;
mem['h0118] = 32'h00D82023;
mem['h0119] = 32'h00052683;
mem['h011A] = 32'h0006A683;
mem['h011B] = 32'h0146A683;
mem['h011C] = 32'h0006A803;
mem['h011D] = 32'h00082683;
mem['h011E] = 32'h0016E693;
mem['h011F] = 32'h00D82023;
mem['h0120] = 32'hF3DFF06F;
mem['h0121] = 32'h00052703;
mem['h0122] = 32'h40D787B3;
mem['h0123] = 32'h000106B7;
mem['h0124] = 32'h00072703;
mem['h0125] = 32'hFFF68693;
mem['h0126] = 32'h40F6D7B3;
mem['h0127] = 32'h01072703;
mem['h0128] = 32'h01079793;
mem['h0129] = 32'h00072603;
mem['h012A] = 32'h00062703;
mem['h012B] = 32'h00D77733;
mem['h012C] = 32'h00F767B3;
mem['h012D] = 32'h00F62023;
mem['h012E] = 32'h00052783;
mem['h012F] = 32'h000086B7;
mem['h0130] = 32'h0007A783;
mem['h0131] = 32'h0107A783;
mem['h0132] = 32'h0007A703;
mem['h0133] = 32'h00072783;
mem['h0134] = 32'h00D7E7B3;
mem['h0135] = 32'h00F72023;
mem['h0136] = 32'h00052783;
mem['h0137] = 32'h0007A783;
mem['h0138] = 32'h0147A783;
mem['h0139] = 32'h0007A703;
mem['h013A] = 32'h00072783;
mem['h013B] = 32'h0017E793;
mem['h013C] = 32'h00F72023;
mem['h013D] = 32'h00008067;
mem['h013E] = 32'hF9010113;
mem['h013F] = 32'h02400513;
mem['h0140] = 32'h06112623;
mem['h0141] = 32'h06812423;
mem['h0142] = 32'h06912223;
mem['h0143] = 32'h07212023;
mem['h0144] = 32'h05312E23;
mem['h0145] = 32'h05412C23;
mem['h0146] = 32'h05512A23;
mem['h0147] = 32'h05612823;
mem['h0148] = 32'h05712623;
mem['h0149] = 32'h05812423;
mem['h014A] = 32'h05912223;
mem['h014B] = 32'h05A12023;
mem['h014C] = 32'h03B12E23;
mem['h014D] = 32'hD59FF0EF;
mem['h014E] = 32'h00050413;
mem['h014F] = 32'h00800513;
mem['h0150] = 32'hD4DFF0EF;
mem['h0151] = 32'h00050913;
mem['h0152] = 32'h01C00513;
mem['h0153] = 32'hD41FF0EF;
mem['h0154] = 32'h00050493;
mem['h0155] = 32'h00400513;
mem['h0156] = 32'hD35FF0EF;
mem['h0157] = 32'h200007B7;
mem['h0158] = 32'h00F52023;
mem['h0159] = 32'h00A4A023;
mem['h015A] = 32'h00400513;
mem['h015B] = 32'hD21FF0EF;
mem['h015C] = 32'h200007B7;
mem['h015D] = 32'h00478793;
mem['h015E] = 32'h00F52023;
mem['h015F] = 32'h00A4A223;
mem['h0160] = 32'h00400513;
mem['h0161] = 32'hD09FF0EF;
mem['h0162] = 32'h200007B7;
mem['h0163] = 32'h00878793;
mem['h0164] = 32'h00F52023;
mem['h0165] = 32'h00A4A423;
mem['h0166] = 32'h00400513;
mem['h0167] = 32'hCF1FF0EF;
mem['h0168] = 32'h200007B7;
mem['h0169] = 32'h00C78793;
mem['h016A] = 32'h00F52023;
mem['h016B] = 32'h00A4A623;
mem['h016C] = 32'h00400513;
mem['h016D] = 32'hCD9FF0EF;
mem['h016E] = 32'h200007B7;
mem['h016F] = 32'h01078793;
mem['h0170] = 32'h00F52023;
mem['h0171] = 32'h00A4A823;
mem['h0172] = 32'h00400513;
mem['h0173] = 32'hCC1FF0EF;
mem['h0174] = 32'h200007B7;
mem['h0175] = 32'h01478793;
mem['h0176] = 32'h00F52023;
mem['h0177] = 32'h00A4AA23;
mem['h0178] = 32'h00400513;
mem['h0179] = 32'hCA9FF0EF;
mem['h017A] = 32'h200007B7;
mem['h017B] = 32'h01878793;
mem['h017C] = 32'h00F52023;
mem['h017D] = 32'h00A4AC23;
mem['h017E] = 32'h00992023;
mem['h017F] = 32'h01C00513;
mem['h0180] = 32'hC8DFF0EF;
mem['h0181] = 32'h00050493;
mem['h0182] = 32'h00400513;
mem['h0183] = 32'hC81FF0EF;
mem['h0184] = 32'h200007B7;
mem['h0185] = 32'h01C78793;
mem['h0186] = 32'h00F52023;
mem['h0187] = 32'h00A4A023;
mem['h0188] = 32'h00400513;
mem['h0189] = 32'hC69FF0EF;
mem['h018A] = 32'h200007B7;
mem['h018B] = 32'h02078793;
mem['h018C] = 32'h00F52023;
mem['h018D] = 32'h00A4A223;
mem['h018E] = 32'h00400513;
mem['h018F] = 32'hC51FF0EF;
mem['h0190] = 32'h200007B7;
mem['h0191] = 32'h02478793;
mem['h0192] = 32'h00F52023;
mem['h0193] = 32'h00A4A423;
mem['h0194] = 32'h00400513;
mem['h0195] = 32'hC39FF0EF;
mem['h0196] = 32'h200007B7;
mem['h0197] = 32'h02878793;
mem['h0198] = 32'h00F52023;
mem['h0199] = 32'h00A4A623;
mem['h019A] = 32'h00400513;
mem['h019B] = 32'hC21FF0EF;
mem['h019C] = 32'h200007B7;
mem['h019D] = 32'h02C78793;
mem['h019E] = 32'h00F52023;
mem['h019F] = 32'h00A4A823;
mem['h01A0] = 32'h00400513;
mem['h01A1] = 32'hC09FF0EF;
mem['h01A2] = 32'h200007B7;
mem['h01A3] = 32'h03078793;
mem['h01A4] = 32'h00F52023;
mem['h01A5] = 32'h00A4AA23;
mem['h01A6] = 32'h00400513;
mem['h01A7] = 32'hBF1FF0EF;
mem['h01A8] = 32'h200007B7;
mem['h01A9] = 32'h03478793;
mem['h01AA] = 32'h00F52023;
mem['h01AB] = 32'h00A4AC23;
mem['h01AC] = 32'h00992223;
mem['h01AD] = 32'h01242023;
mem['h01AE] = 32'h01000513;
mem['h01AF] = 32'hBD1FF0EF;
mem['h01B0] = 32'h00050493;
mem['h01B1] = 32'h00400513;
mem['h01B2] = 32'hBC5FF0EF;
mem['h01B3] = 32'h200007B7;
mem['h01B4] = 32'h03878793;
mem['h01B5] = 32'h00F52023;
mem['h01B6] = 32'h00A4A023;
mem['h01B7] = 32'h00400513;
mem['h01B8] = 32'hBADFF0EF;
mem['h01B9] = 32'h200007B7;
mem['h01BA] = 32'h03C78793;
mem['h01BB] = 32'h00F52023;
mem['h01BC] = 32'h00A4A223;
mem['h01BD] = 32'h00400513;
mem['h01BE] = 32'hB95FF0EF;
mem['h01BF] = 32'h200007B7;
mem['h01C0] = 32'h04078793;
mem['h01C1] = 32'h00F52023;
mem['h01C2] = 32'h00A4A423;
mem['h01C3] = 32'h00400513;
mem['h01C4] = 32'hB7DFF0EF;
mem['h01C5] = 32'h200007B7;
mem['h01C6] = 32'h04478793;
mem['h01C7] = 32'h00F52023;
mem['h01C8] = 32'h00A4A623;
mem['h01C9] = 32'h00942223;
mem['h01CA] = 32'h00400513;
mem['h01CB] = 32'hB61FF0EF;
mem['h01CC] = 32'h200007B7;
mem['h01CD] = 32'h04878793;
mem['h01CE] = 32'h00F52023;
mem['h01CF] = 32'h200004B7;
mem['h01D0] = 32'hE0000A37;
mem['h01D1] = 32'h200009B7;
mem['h01D2] = 32'h00A42423;
mem['h01D3] = 32'h04C48493;
mem['h01D4] = 32'hFC0A0A13;
mem['h01D5] = 32'h05C98993;
mem['h01D6] = 32'h00400513;
mem['h01D7] = 32'hB31FF0EF;
mem['h01D8] = 32'h00050913;
mem['h01D9] = 32'h00400513;
mem['h01DA] = 32'hB25FF0EF;
mem['h01DB] = 32'h00952023;
mem['h01DC] = 32'h014487B3;
mem['h01DD] = 32'h00A92023;
mem['h01DE] = 32'h00F407B3;
mem['h01DF] = 32'h0127A023;
mem['h01E0] = 32'h00448493;
mem['h01E1] = 32'hFD349AE3;
mem['h01E2] = 32'h00400513;
mem['h01E3] = 32'hB01FF0EF;
mem['h01E4] = 32'h00050913;
mem['h01E5] = 32'h00400513;
mem['h01E6] = 32'hAF5FF0EF;
mem['h01E7] = 32'h00952023;
mem['h01E8] = 32'h00A92023;
mem['h01E9] = 32'h01242E23;
mem['h01EA] = 32'h00400513;
mem['h01EB] = 32'hAE1FF0EF;
mem['h01EC] = 32'h200007B7;
mem['h01ED] = 32'h06078793;
mem['h01EE] = 32'h00F52023;
mem['h01EF] = 32'h000014B7;
mem['h01F0] = 32'hEFC48593;
mem['h01F1] = 32'h02A42023;
mem['h01F2] = 32'h00040513;
mem['h01F3] = 32'hA05FF0EF;
mem['h01F4] = 32'h000015B7;
mem['h01F5] = 32'hF2C58593;
mem['h01F6] = 32'h00040513;
mem['h01F7] = 32'h9F5FF0EF;
mem['h01F8] = 32'hEFC48593;
mem['h01F9] = 32'h00040513;
mem['h01FA] = 32'h9E9FF0EF;
mem['h01FB] = 32'h000015B7;
mem['h01FC] = 32'hF5C58593;
mem['h01FD] = 32'h00040513;
mem['h01FE] = 32'h9D9FF0EF;
mem['h01FF] = 32'h000015B7;
mem['h0200] = 32'hF7458593;
mem['h0201] = 32'h00040513;
mem['h0202] = 32'h9C9FF0EF;
mem['h0203] = 32'h10000937;
mem['h0204] = 32'h00090593;
mem['h0205] = 32'h00040513;
mem['h0206] = 32'h9FDFF0EF;
mem['h0207] = 32'h000015B7;
mem['h0208] = 32'hF8C58593;
mem['h0209] = 32'h00040513;
mem['h020A] = 32'h00090493;
mem['h020B] = 32'h9A5FF0EF;
mem['h020C] = 32'h00448593;
mem['h020D] = 32'h00040513;
mem['h020E] = 32'h9DDFF0EF;
mem['h020F] = 32'h000015B7;
mem['h0210] = 32'hFA858593;
mem['h0211] = 32'h00040513;
mem['h0212] = 32'h989FF0EF;
mem['h0213] = 32'h0084C583;
mem['h0214] = 32'h00200613;
mem['h0215] = 32'h00040513;
mem['h0216] = 32'h845FF0EF;
mem['h0217] = 32'h03A00593;
mem['h0218] = 32'h00040513;
mem['h0219] = 32'h811FF0EF;
mem['h021A] = 32'h0094C583;
mem['h021B] = 32'h00200613;
mem['h021C] = 32'h00040513;
mem['h021D] = 32'h829FF0EF;
mem['h021E] = 32'h03A00593;
mem['h021F] = 32'h00040513;
mem['h0220] = 32'hFF4FF0EF;
mem['h0221] = 32'h00A4C583;
mem['h0222] = 32'h00200613;
mem['h0223] = 32'h00040513;
mem['h0224] = 32'h80DFF0EF;
mem['h0225] = 32'h03A00593;
mem['h0226] = 32'h00040513;
mem['h0227] = 32'hFD8FF0EF;
mem['h0228] = 32'h00B4C583;
mem['h0229] = 32'h00200613;
mem['h022A] = 32'h00040513;
mem['h022B] = 32'hFF0FF0EF;
mem['h022C] = 32'h03A00593;
mem['h022D] = 32'h00040513;
mem['h022E] = 32'hFBCFF0EF;
mem['h022F] = 32'h00C4C583;
mem['h0230] = 32'h00200613;
mem['h0231] = 32'h00040513;
mem['h0232] = 32'hFD4FF0EF;
mem['h0233] = 32'h03A00593;
mem['h0234] = 32'h00040513;
mem['h0235] = 32'hFA0FF0EF;
mem['h0236] = 32'h00D4C583;
mem['h0237] = 32'h00200613;
mem['h0238] = 32'h00040513;
mem['h0239] = 32'hFB8FF0EF;
mem['h023A] = 32'h000015B7;
mem['h023B] = 32'hFC458593;
mem['h023C] = 32'h00040513;
mem['h023D] = 32'h8DDFF0EF;
mem['h023E] = 32'h00E48593;
mem['h023F] = 32'h00040513;
mem['h0240] = 32'h915FF0EF;
mem['h0241] = 32'h000015B7;
mem['h0242] = 32'hFE058593;
mem['h0243] = 32'h00040513;
mem['h0244] = 32'h8C1FF0EF;
mem['h0245] = 32'h0124C583;
mem['h0246] = 32'h00040513;
mem['h0247] = 32'h000014B7;
mem['h0248] = 32'hFE8FF0EF;
mem['h0249] = 32'hFFC48593;
mem['h024A] = 32'h00040513;
mem['h024B] = 32'h8A5FF0EF;
mem['h024C] = 32'h000015B7;
mem['h024D] = 32'h00058593;
mem['h024E] = 32'h00040513;
mem['h024F] = 32'h100009B7;
mem['h0250] = 32'h891FF0EF;
mem['h0251] = 32'h01898B93;
mem['h0252] = 32'h608B8793;
mem['h0253] = 32'h00090A13;
mem['h0254] = 32'h00F12623;
mem['h0255] = 32'h00A00A93;
mem['h0256] = 32'h00D00B13;
mem['h0257] = 32'h000B8023;
mem['h0258] = 32'h000B9123;
mem['h0259] = 32'h00042703;
mem['h025A] = 32'h00472703;
mem['h025B] = 32'h01872703;
mem['h025C] = 32'h00072703;
mem['h025D] = 32'h00072703;
mem['h025E] = 32'h00177713;
mem['h025F] = 32'h0E070863;
mem['h0260] = 32'h00042703;
mem['h0261] = 32'h000B8C93;
mem['h0262] = 32'h01898693;
mem['h0263] = 32'h00472703;
mem['h0264] = 32'h01072703;
mem['h0265] = 32'h00072703;
mem['h0266] = 32'h00072703;
mem['h0267] = 32'h00375713;
mem['h0268] = 32'h00777713;
mem['h0269] = 32'h00EB80A3;
mem['h026A] = 32'h00000713;
mem['h026B] = 32'h00042603;
mem['h026C] = 32'h01068693;
mem['h026D] = 32'h00462603;
mem['h026E] = 32'h00062603;
mem['h026F] = 32'h00062603;
mem['h0270] = 32'h00062603;
mem['h0271] = 32'hFEC6AC23;
mem['h0272] = 32'h00042603;
mem['h0273] = 32'h00462603;
mem['h0274] = 32'h00462603;
mem['h0275] = 32'h00062603;
mem['h0276] = 32'h00062603;
mem['h0277] = 32'hFEC6AE23;
mem['h0278] = 32'h00042603;
mem['h0279] = 32'h00462603;
mem['h027A] = 32'h00862603;
mem['h027B] = 32'h00062603;
mem['h027C] = 32'h00062603;
mem['h027D] = 32'h00C6A023;
mem['h027E] = 32'h00042603;
mem['h027F] = 32'h00462603;
mem['h0280] = 32'h00C62603;
mem['h0281] = 32'h00062603;
mem['h0282] = 32'h00062603;
mem['h0283] = 32'h00C6A223;
mem['h0284] = 32'h00042603;
mem['h0285] = 32'h00462603;
mem['h0286] = 32'h01062603;
mem['h0287] = 32'h00062603;
mem['h0288] = 32'h00062603;
mem['h0289] = 32'h01061593;
mem['h028A] = 32'h0605D463;
mem['h028B] = 32'h00042683;
mem['h028C] = 32'h0046A683;
mem['h028D] = 32'h0106A683;
mem['h028E] = 32'h0006A683;
mem['h028F] = 32'h0026D683;
mem['h0290] = 32'h0016F613;
mem['h0291] = 32'h04061063;
mem['h0292] = 32'h00042683;
mem['h0293] = 32'h00EBA223;
mem['h0294] = 32'h0046A683;
mem['h0295] = 32'h0146A683;
mem['h0296] = 32'h0006A603;
mem['h0297] = 32'h00062683;
mem['h0298] = 32'h0016E693;
mem['h0299] = 32'h00D62023;
mem['h029A] = 32'h04071663;
mem['h029B] = 32'h00842703;
mem['h029C] = 32'h00072683;
mem['h029D] = 32'h0006A703;
mem['h029E] = 32'hDFF77713;
mem['h029F] = 32'h00E6A023;
mem['h02A0] = 32'h0D00006F;
mem['h02A1] = 32'h00170713;
mem['h02A2] = 32'h0016D693;
mem['h02A3] = 32'hFB5FF06F;
mem['h02A4] = 32'h00042603;
mem['h02A5] = 32'h01070713;
mem['h02A6] = 32'h00462603;
mem['h02A7] = 32'h01462603;
mem['h02A8] = 32'h00062583;
mem['h02A9] = 32'h0005A603;
mem['h02AA] = 32'h00166613;
mem['h02AB] = 32'h00C5A023;
mem['h02AC] = 32'hEFDFF06F;
mem['h02AD] = 32'h00842703;
mem['h02AE] = 32'h00072683;
mem['h02AF] = 32'h0006A703;
mem['h02B0] = 32'h20076713;
mem['h02B1] = 32'h00E6A023;
mem['h02B2] = 32'h014BCD03;
mem['h02B3] = 32'h00800713;
mem['h02B4] = 32'h04ED1E63;
mem['h02B5] = 32'h015BC703;
mem['h02B6] = 32'h00600693;
mem['h02B7] = 32'h0AD70463;
mem['h02B8] = 32'h04071663;
mem['h02B9] = 32'h016BC703;
mem['h02BA] = 32'h04000693;
mem['h02BB] = 32'h0F077713;
mem['h02BC] = 32'h02D71E63;
mem['h02BD] = 32'h01FBC683;
mem['h02BE] = 32'h00100713;
mem['h02BF] = 32'h02E69863;
mem['h02C0] = 32'h000017B7;
mem['h02C1] = 32'h03078593;
mem['h02C2] = 32'h00040513;
mem['h02C3] = 32'hEC4FF0EF;
mem['h02C4] = 32'h004BA583;
mem['h02C5] = 32'h00400613;
mem['h02C6] = 32'h00040513;
mem['h02C7] = 32'hD80FF0EF;
mem['h02C8] = 32'hFFC48593;
mem['h02C9] = 32'h00040513;
mem['h02CA] = 32'hEA8FF0EF;
mem['h02CB] = 32'h001BC683;
mem['h02CC] = 32'h00100713;
mem['h02CD] = 32'h1AE69463;
mem['h02CE] = 32'h00200713;
mem['h02CF] = 32'h00EB8023;
mem['h02D0] = 32'h00DB81A3;
mem['h02D1] = 32'h01898593;
mem['h02D2] = 32'h00040513;
mem['h02D3] = 32'hF94FF0EF;
mem['h02D4] = 32'h00442703;
mem['h02D5] = 32'h00072703;
mem['h02D6] = 32'h00072703;
mem['h02D7] = 32'h00072583;
mem['h02D8] = 32'hDE05DEE3;
mem['h02D9] = 32'h0FF5F713;
mem['h02DA] = 32'h01200693;
mem['h02DB] = 32'hDED708E3;
mem['h02DC] = 32'h0FF5F593;
mem['h02DD] = 32'h00B10823;
mem['h02DE] = 32'h17559C63;
mem['h02DF] = 32'h00010823;
mem['h02E0] = 32'hDDDFF06F;
mem['h02E1] = 32'h000017B7;
mem['h02E2] = 32'h04478593;
mem['h02E3] = 32'h00040513;
mem['h02E4] = 32'hE40FF0EF;
mem['h02E5] = 32'h004BC583;
mem['h02E6] = 32'h00040513;
mem['h02E7] = 32'hD6CFF0EF;
mem['h02E8] = 32'hFFC48593;
mem['h02E9] = 32'h00040513;
mem['h02EA] = 32'hE28FF0EF;
mem['h02EB] = 32'h017BC683;
mem['h02EC] = 32'h00100613;
mem['h02ED] = 32'h016BC703;
mem['h02EE] = 32'hF6C69AE3;
mem['h02EF] = 32'h018BC603;
mem['h02F0] = 32'hF7A616E3;
mem['h02F1] = 32'h019BC603;
mem['h02F2] = 32'h00C76733;
mem['h02F3] = 32'h01CBC603;
mem['h02F4] = 32'h00C76733;
mem['h02F5] = 32'hF4071CE3;
mem['h02F6] = 32'h01DBC703;
mem['h02F7] = 32'hF4D718E3;
mem['h02F8] = 32'h00000693;
mem['h02F9] = 32'h00400593;
mem['h02FA] = 32'h00DA0633;
mem['h02FB] = 32'h02ECC703;
mem['h02FC] = 32'h00064603;
mem['h02FD] = 32'h0CC70A63;
mem['h02FE] = 32'h40C70733;
mem['h02FF] = 32'h001BC683;
mem['h0300] = 32'hF20716E3;
mem['h0301] = 32'h00100713;
mem['h0302] = 32'h60EB85A3;
mem['h0303] = 32'h81E18593;
mem['h0304] = 32'h02A00713;
mem['h0305] = 32'h610B8513;
mem['h0306] = 32'h00600613;
mem['h0307] = 32'h60DB8423;
mem['h0308] = 32'h60EBA623;
mem['h0309] = 32'hE9CFF0EF;
mem['h030A] = 32'h008A0593;
mem['h030B] = 32'h616B8513;
mem['h030C] = 32'h00600613;
mem['h030D] = 32'hE8CFF0EF;
mem['h030E] = 32'h01000737;
mem['h030F] = 32'h60870713;
mem['h0310] = 32'h60EBAE23;
mem['h0311] = 32'h04060737;
mem['h0312] = 32'h100007B7;
mem['h0313] = 32'h00870713;
mem['h0314] = 32'h00878593;
mem['h0315] = 32'h62EBA023;
mem['h0316] = 32'h626B8513;
mem['h0317] = 32'h20000713;
mem['h0318] = 32'h00600613;
mem['h0319] = 32'h62EB9223;
mem['h031A] = 32'hE58FF0EF;
mem['h031B] = 32'h00090593;
mem['h031C] = 32'h62CB8513;
mem['h031D] = 32'h00400613;
mem['h031E] = 32'hE48FF0EF;
mem['h031F] = 32'h81E18593;
mem['h0320] = 32'h630B8513;
mem['h0321] = 32'h00600613;
mem['h0322] = 32'hE38FF0EF;
mem['h0323] = 32'h00400613;
mem['h0324] = 32'h024B8593;
mem['h0325] = 32'h636B8513;
mem['h0326] = 32'hE28FF0EF;
mem['h0327] = 32'h00C12583;
mem['h0328] = 32'h00040513;
mem['h0329] = 32'hE3CFF0EF;
mem['h032A] = 32'h000017B7;
mem['h032B] = 32'h05878593;
mem['h032C] = 32'h00040513;
mem['h032D] = 32'hD1CFF0EF;
mem['h032E] = 32'h60CBC583;
mem['h032F] = 32'h00040513;
mem['h0330] = 32'hC48FF0EF;
mem['h0331] = 32'hE5DFF06F;
mem['h0332] = 32'h00168693;
mem['h0333] = 32'h001C8C93;
mem['h0334] = 32'hF0B69CE3;
mem['h0335] = 32'h00000713;
mem['h0336] = 32'hF25FF06F;
mem['h0337] = 32'h00200613;
mem['h0338] = 32'hE6C698E3;
mem['h0339] = 32'h00EB8023;
mem['h033A] = 32'h00EB81A3;
mem['h033B] = 32'hE59FF06F;
mem['h033C] = 32'h00000C93;
mem['h033D] = 32'h01010C13;
mem['h033E] = 32'h07658863;
mem['h033F] = 32'h00800D13;
mem['h0340] = 32'h07F00D93;
mem['h0341] = 32'h01A58463;
mem['h0342] = 32'h0FB59A63;
mem['h0343] = 32'h03905863;
mem['h0344] = 32'h00800593;
mem['h0345] = 32'h00040513;
mem['h0346] = 32'hB5CFF0EF;
mem['h0347] = 32'h02000593;
mem['h0348] = 32'h00040513;
mem['h0349] = 32'hB50FF0EF;
mem['h034A] = 32'h00800593;
mem['h034B] = 32'h00040513;
mem['h034C] = 32'hFFFC0C13;
mem['h034D] = 32'hFFFC8C93;
mem['h034E] = 32'hB3CFF0EF;
mem['h034F] = 32'h00442603;
mem['h0350] = 32'h00062603;
mem['h0351] = 32'h00062603;
mem['h0352] = 32'h00062583;
mem['h0353] = 32'hFE05D8E3;
mem['h0354] = 32'h01F00793;
mem['h0355] = 32'h02FC8663;
mem['h0356] = 32'h0FF5F593;
mem['h0357] = 32'h00BC0023;
mem['h0358] = 32'h03558063;
mem['h0359] = 32'hFB6590E3;
mem['h035A] = 32'h00D00593;
mem['h035B] = 32'h00040513;
mem['h035C] = 32'hB04FF0EF;
mem['h035D] = 32'h00A00593;
mem['h035E] = 32'h00040513;
mem['h035F] = 32'hAF8FF0EF;
mem['h0360] = 32'h000C0023;
mem['h0361] = 32'h0FFCFC93;
mem['h0362] = 32'hBC0C8AE3;
mem['h0363] = 32'h000015B7;
mem['h0364] = 32'h00040513;
mem['h0365] = 32'h06C58593;
mem['h0366] = 32'hC38FF0EF;
mem['h0367] = 32'h01010593;
mem['h0368] = 32'h00040513;
mem['h0369] = 32'hC2CFF0EF;
mem['h036A] = 32'hFFC48593;
mem['h036B] = 32'h00040513;
mem['h036C] = 32'hC20FF0EF;
mem['h036D] = 32'h000015B7;
mem['h036E] = 32'h00040513;
mem['h036F] = 32'h07858593;
mem['h0370] = 32'hC10FF0EF;
mem['h0371] = 32'h000C8593;
mem['h0372] = 32'h00040513;
mem['h0373] = 32'hB3CFF0EF;
mem['h0374] = 32'hFFC48593;
mem['h0375] = 32'h00040513;
mem['h0376] = 32'hBF8FF0EF;
mem['h0377] = 32'h01014583;
mem['h0378] = 32'h00040513;
mem['h0379] = 32'h00200613;
mem['h037A] = 32'hAB4FF0EF;
mem['h037B] = 32'hFFC48593;
mem['h037C] = 32'h00040513;
mem['h037D] = 32'hBDCFF0EF;
mem['h037E] = 32'hB5DFF06F;
mem['h037F] = 32'h00040513;
mem['h0380] = 32'hA74FF0EF;
mem['h0381] = 32'h001C0C13;
mem['h0382] = 32'h001C8C93;
mem['h0383] = 32'hF31FF06F;
mem['h0384] = 32'h00050613;
mem['h0385] = 32'h00000513;
mem['h0386] = 32'h0015F693;
mem['h0387] = 32'h00068463;
mem['h0388] = 32'h00C50533;
mem['h0389] = 32'h0015D593;
mem['h038A] = 32'h00161613;
mem['h038B] = 32'hFE0596E3;
mem['h038C] = 32'h00008067;
mem['h038D] = 32'h06054063;
mem['h038E] = 32'h0605C663;
mem['h038F] = 32'h00058613;
mem['h0390] = 32'h00050593;
mem['h0391] = 32'hFFF00513;
mem['h0392] = 32'h02060C63;
mem['h0393] = 32'h00100693;
mem['h0394] = 32'h00B67A63;
mem['h0395] = 32'h00C05863;
mem['h0396] = 32'h00161613;
mem['h0397] = 32'h00169693;
mem['h0398] = 32'hFEB66AE3;
mem['h0399] = 32'h00000513;
mem['h039A] = 32'h00C5E663;
mem['h039B] = 32'h40C585B3;
mem['h039C] = 32'h00D56533;
mem['h039D] = 32'h0016D693;
mem['h039E] = 32'h00165613;
mem['h039F] = 32'hFE0696E3;
mem['h03A0] = 32'h00008067;
mem['h03A1] = 32'h00008293;
mem['h03A2] = 32'hFB5FF0EF;
mem['h03A3] = 32'h00058513;
mem['h03A4] = 32'h00028067;
mem['h03A5] = 32'h40A00533;
mem['h03A6] = 32'h00B04863;
mem['h03A7] = 32'h40B005B3;
mem['h03A8] = 32'hF9DFF06F;
mem['h03A9] = 32'h40B005B3;
mem['h03AA] = 32'h00008293;
mem['h03AB] = 32'hF91FF0EF;
mem['h03AC] = 32'h40A00533;
mem['h03AD] = 32'h00028067;
mem['h03AE] = 32'h00008293;
mem['h03AF] = 32'h0005CA63;
mem['h03B0] = 32'h00054C63;
mem['h03B1] = 32'hF79FF0EF;
mem['h03B2] = 32'h00058513;
mem['h03B3] = 32'h00028067;
mem['h03B4] = 32'h40B005B3;
mem['h03B5] = 32'hFE0558E3;
mem['h03B6] = 32'h40A00533;
mem['h03B7] = 32'hF61FF0EF;
mem['h03B8] = 32'h40B00533;
mem['h03B9] = 32'h00028067;
mem['h03BA] = 32'h33323130;
mem['h03BB] = 32'h37363534;
mem['h03BC] = 32'h42413938;
mem['h03BD] = 32'h46454443;
mem['h03BE] = 32'h00000000;
mem['h03BF] = 32'h3D3D3D3D;
mem['h03C0] = 32'h3D3D3D3D;
mem['h03C1] = 32'h3D3D3D3D;
mem['h03C2] = 32'h3D3D3D3D;
mem['h03C3] = 32'h3D3D3D3D;
mem['h03C4] = 32'h3D3D3D3D;
mem['h03C5] = 32'h3D3D3D3D;
mem['h03C6] = 32'h3D3D3D3D;
mem['h03C7] = 32'h3D3D3D3D;
mem['h03C8] = 32'h3D3D3D3D;
mem['h03C9] = 32'h0A0D3D3D;
mem['h03CA] = 32'h00000000;
mem['h03CB] = 32'h20202020;
mem['h03CC] = 32'h57202020;
mem['h03CD] = 32'h47657269;
mem['h03CE] = 32'h64726175;
mem['h03CF] = 32'h47504620;
mem['h03D0] = 32'h79622041;
mem['h03D1] = 32'h69684320;
mem['h03D2] = 32'h6843696C;
mem['h03D3] = 32'h20737069;
mem['h03D4] = 32'h20202020;
mem['h03D5] = 32'h0A0D2020;
mem['h03D6] = 32'h00000000;
mem['h03D7] = 32'h7774654E;
mem['h03D8] = 32'h206B726F;
mem['h03D9] = 32'h666E6F63;
mem['h03DA] = 32'h72756769;
mem['h03DB] = 32'h6F697461;
mem['h03DC] = 32'h000A0D6E;
mem['h03DD] = 32'h49202D2D;
mem['h03DE] = 32'h64612050;
mem['h03DF] = 32'h73657264;
mem['h03E0] = 32'h20203A73;
mem['h03E1] = 32'h20202020;
mem['h03E2] = 32'h00002020;
mem['h03E3] = 32'h2D2D0A0D;
mem['h03E4] = 32'h62755320;
mem['h03E5] = 32'h2074656E;
mem['h03E6] = 32'h6B73616D;
mem['h03E7] = 32'h2020203A;
mem['h03E8] = 32'h20202020;
mem['h03E9] = 32'h00000000;
mem['h03EA] = 32'h2D2D0A0D;
mem['h03EB] = 32'h43414D20;
mem['h03EC] = 32'h64646120;
mem['h03ED] = 32'h73736572;
mem['h03EE] = 32'h2020203A;
mem['h03EF] = 32'h20202020;
mem['h03F0] = 32'h00000000;
mem['h03F1] = 32'h2D2D0A0D;
mem['h03F2] = 32'h66654420;
mem['h03F3] = 32'h746C7561;
mem['h03F4] = 32'h74616720;
mem['h03F5] = 32'h79617765;
mem['h03F6] = 32'h2020203A;
mem['h03F7] = 32'h00000000;
mem['h03F8] = 32'h2D2D0A0D;
mem['h03F9] = 32'h66654420;
mem['h03FA] = 32'h746C7561;
mem['h03FB] = 32'h746E6920;
mem['h03FC] = 32'h61667265;
mem['h03FD] = 32'h203A6563;
mem['h03FE] = 32'h00000000;
mem['h03FF] = 32'h00000A0D;
mem['h0400] = 32'h2D2D2D2D;
mem['h0401] = 32'h2D2D2D2D;
mem['h0402] = 32'h2D2D2D2D;
mem['h0403] = 32'h2D2D2D2D;
mem['h0404] = 32'h2D2D2D2D;
mem['h0405] = 32'h2D2D2D2D;
mem['h0406] = 32'h2D2D2D2D;
mem['h0407] = 32'h2D2D2D2D;
mem['h0408] = 32'h2D2D2D2D;
mem['h0409] = 32'h2D2D2D2D;
mem['h040A] = 32'h0A0D2D2D;
mem['h040B] = 32'h00000000;
mem['h040C] = 32'h5F54454E;
mem['h040D] = 32'h544F5250;
mem['h040E] = 32'h43495F4F;
mem['h040F] = 32'h203A504D;
mem['h0410] = 32'h00000000;
mem['h0411] = 32'h4E203C3C;
mem['h0412] = 32'h505F5445;
mem['h0413] = 32'h4F544F52;
mem['h0414] = 32'h5052415F;
mem['h0415] = 32'h0000203A;
mem['h0416] = 32'h4E203E3E;
mem['h0417] = 32'h505F5445;
mem['h0418] = 32'h4F544F52;
mem['h0419] = 32'h5052415F;
mem['h041A] = 32'h0000203A;
mem['h041B] = 32'h65636552;
mem['h041C] = 32'h64657669;
mem['h041D] = 32'h0000203A;
mem['h041E] = 32'h65636552;
mem['h041F] = 32'h64657669;
mem['h0420] = 32'h6E656C20;
mem['h0421] = 32'h3A687467;
mem['h0422] = 32'h00000020;
mem['h0423] = 32'h6301A8C0;
mem['h0424] = 32'h00FFFFFF;
mem['h0425] = 32'hAECCCACA;
mem['h0426] = 32'hA8C00100;
mem['h0427] = 32'h0001FE01;
mem['h0428] = 32'h00000000;
