-- Timing params:
--   Fixed?: False
--   Pipeline Slices: [0.07692307692307693, 0.15384615384615385, 0.23076923076923078, 0.3076923076923077, 0.38461538461538464, 0.46153846153846156, 0.5384615384615385, 0.6153846153846154, 0.6923076923076923, 0.7692307692307692, 0.846153846153846, 0.9230769230769229]
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 3
entity chacha20_decrypt_pipeline_no_handshake_12CLK_e61aba39 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 global_to_module : in chacha20_decrypt_pipeline_no_handshake_global_to_module_t;
 module_to_global : out chacha20_decrypt_pipeline_no_handshake_module_to_global_t);
end chacha20_decrypt_pipeline_no_handshake_12CLK_e61aba39;
architecture arch of chacha20_decrypt_pipeline_no_handshake_12CLK_e61aba39 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 12;
-- All of the wires/regs in function
-- Stage 0
signal REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 1
signal REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 2
signal REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 3
signal REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 4
signal REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 5
signal REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 6
signal REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 7
signal REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 8
signal REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 9
signal REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 10
signal REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Stage 11
signal REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- chacha20_decrypt_pipeline_no_handshake_in_reg_func[chacha20_decrypt_c_l24_c102_ef13]
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_CLOCK_ENABLE : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_data : chacha20_decrypt_loop_body_in_t;
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_id : unsigned(7 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_valid : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output : chacha20_decrypt_pipeline_no_handshake_in_reg_t;

-- chacha20_decrypt_loop_body[chacha20_decrypt_c_l24_c308_fc66]
signal chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_inputs : chacha20_decrypt_loop_body_in_t;
signal chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output : axis512_t;

-- chacha20_decrypt_pipeline_no_handshake_out_reg_func[chacha20_decrypt_c_l24_c397_ca6f]
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_data : axis512_t;
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
signal chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output : chacha20_decrypt_pipeline_no_handshake_out_reg_t;


begin

-- SUBMODULE INSTANCES 
-- chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13 : 0 clocks latency
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13 : entity work.chacha20_decrypt_pipeline_no_handshake_in_reg_func_0CLK_b45f1687 port map (
clk,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_CLOCK_ENABLE,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_data,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_id,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_valid,
chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output);

-- chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66 : 12 clocks latency
chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66 : entity work.chacha20_decrypt_loop_body_12CLK_e38dbbb7 port map (
clk,
chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_inputs,
chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output);

-- chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f : 0 clocks latency
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f : entity work.chacha20_decrypt_pipeline_no_handshake_out_reg_func_0CLK_b45f1687 port map (
clk,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_data,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Registers
 -- Stage 0
 REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 1
 REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 2
 REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 3
 REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 4
 REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 5
 REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 6
 REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 7
 REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 8
 REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 9
 REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 10
 REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Stage 11
 REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id,
 REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid,
 REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE,
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output,
 chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output,
 chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in : chacha20_decrypt_loop_body_in_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_valid : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out : axis512_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_valid : unsigned(0 downto 0);
 variable VAR_i : chacha20_decrypt_pipeline_no_handshake_in_reg_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_data : chacha20_decrypt_loop_body_in_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_valid : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output : chacha20_decrypt_pipeline_no_handshake_in_reg_t;
 variable VAR_d : axis512_t;
 variable VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_inputs : chacha20_decrypt_loop_body_in_t;
 variable VAR_CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d_chacha20_decrypt_c_l24_c335_2fb4_return_output : chacha20_decrypt_loop_body_in_t;
 variable VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output : axis512_t;
 variable VAR_o : chacha20_decrypt_pipeline_no_handshake_out_reg_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_data : axis512_t;
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id : unsigned(7 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d_chacha20_decrypt_c_l24_c453_eb25_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d_chacha20_decrypt_c_l24_c459_c772_return_output : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output : chacha20_decrypt_pipeline_no_handshake_out_reg_t;
 variable VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d_chacha20_decrypt_c_l24_c515_9c10_return_output : axis512_t;
 variable VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d_chacha20_decrypt_c_l24_c571_01eb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d_chacha20_decrypt_c_l24_c628_4124_return_output : unsigned(0 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_id := to_unsigned(0, 8);
 -- Reads from global variables
     VAR_chacha20_decrypt_pipeline_no_handshake_in := global_to_module.chacha20_decrypt_pipeline_no_handshake_in;
     VAR_chacha20_decrypt_pipeline_no_handshake_in_valid := global_to_module.chacha20_decrypt_pipeline_no_handshake_in_valid;
     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_valid := VAR_chacha20_decrypt_pipeline_no_handshake_in_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_data := VAR_chacha20_decrypt_pipeline_no_handshake_in;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;

     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := VAR_CLOCK_ENABLE;
     -- chacha20_decrypt_pipeline_no_handshake_in_reg_func[chacha20_decrypt_c_l24_c102_ef13] LATENCY=0
     -- Clock enable
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_CLOCK_ENABLE;
     -- Inputs
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_data <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_data;
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_id <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_id;
     chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_valid;
     -- Outputs
     VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output := chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output;

     -- Submodule level 1
     -- CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d[chacha20_decrypt_c_l24_c453_eb25] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d_chacha20_decrypt_c_l24_c453_eb25_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output.id;

     -- CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d[chacha20_decrypt_c_l24_c459_c772] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d_chacha20_decrypt_c_l24_c459_c772_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output.valid;

     -- CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d[chacha20_decrypt_c_l24_c335_2fb4] LATENCY=0
     VAR_CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d_chacha20_decrypt_c_l24_c335_2fb4_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_in_reg_func_chacha20_decrypt_c_l24_c102_ef13_return_output.data;

     -- Submodule level 2
     VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_inputs := VAR_CONST_REF_RD_chacha20_decrypt_loop_body_in_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_data_d41d_chacha20_decrypt_c_l24_c335_2fb4_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_valid_d41d_chacha20_decrypt_c_l24_c459_c772_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_in_reg_t_id_d41d_chacha20_decrypt_c_l24_c453_eb25_return_output;
     -- chacha20_decrypt_loop_body[chacha20_decrypt_c_l24_c308_fc66] LATENCY=12
     -- Inputs
     chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_inputs <= VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_inputs;

     -- Write to comb signals
     COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 1 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 2 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 3 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 4 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 5 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 6 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 7 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 8 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 9 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 10 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 11 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;

     -- Write to comb signals
     COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
   elsif STAGE = 12 then
     -- Read from prev stage
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id := REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid := REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE := REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Submodule outputs
     VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output := chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output;

     -- Submodule level 0
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_data := VAR_chacha20_decrypt_loop_body_chacha20_decrypt_c_l24_c308_fc66_return_output;
     -- chacha20_decrypt_pipeline_no_handshake_out_reg_func[chacha20_decrypt_c_l24_c397_ca6f] LATENCY=0
     -- Clock enable
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Inputs
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_data <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_data;
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     -- Outputs
     VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output := chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output;

     -- Submodule level 1
     -- CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d[chacha20_decrypt_c_l24_c515_9c10] LATENCY=0
     VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d_chacha20_decrypt_c_l24_c515_9c10_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output.data;

     -- CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d[chacha20_decrypt_c_l24_c628_4124] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d_chacha20_decrypt_c_l24_c628_4124_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output.valid;

     -- CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d[chacha20_decrypt_c_l24_c571_01eb] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d_chacha20_decrypt_c_l24_c571_01eb_return_output := VAR_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_return_output.id;

     -- Submodule level 2
     VAR_chacha20_decrypt_pipeline_no_handshake_out := VAR_CONST_REF_RD_axis512_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_data_d41d_chacha20_decrypt_c_l24_c515_9c10_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_valid := VAR_CONST_REF_RD_uint1_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_valid_d41d_chacha20_decrypt_c_l24_c628_4124_return_output;
     VAR_chacha20_decrypt_pipeline_no_handshake_out_id := VAR_CONST_REF_RD_uint8_t_chacha20_decrypt_pipeline_no_handshake_out_reg_t_id_d41d_chacha20_decrypt_c_l24_c571_01eb_return_output;
   end if;
 end loop;

-- Global wires driven various places in pipeline
if clk_en_internal='1' then
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out <= VAR_chacha20_decrypt_pipeline_no_handshake_out;
else
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out <= axis512_t_NULL;
end if;
if clk_en_internal='1' then
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out_valid <= VAR_chacha20_decrypt_pipeline_no_handshake_out_valid;
else
  module_to_global.chacha20_decrypt_pipeline_no_handshake_out_valid <= to_unsigned(0, 1);
end if;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     -- Stage 0
     REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE0_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 1
     REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE1_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 2
     REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE2_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 3
     REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE3_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 4
     REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE4_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 5
     REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE5_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 6
     REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE6_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 7
     REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE7_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 8
     REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE8_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 9
     REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE9_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 10
     REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE10_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
     -- Stage 11
     REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id <= COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_id;
     REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid <= COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_valid;
     REG_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE <= COMB_STAGE11_chacha20_decrypt_pipeline_no_handshake_out_reg_func_chacha20_decrypt_c_l24_c397_ca6f_CLOCK_ENABLE;
 end if;
 end if;
end process;

end arch;
