mem['h0000] = 32'h00000517;
mem['h0001] = 32'h3FC50513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h00418593;
mem['h000F] = 32'h00B55863;
mem['h0010] = 32'h00052023;
mem['h0011] = 32'h00450513;
mem['h0012] = 32'hFEB54CE3;
mem['h0013] = 32'h10008117;
mem['h0014] = 32'hFB410113;
mem['h0015] = 32'h10000197;
mem['h0016] = 32'h7AC18193;
mem['h0017] = 32'h00A54533;
mem['h0018] = 32'h00B5C5B3;
mem['h0019] = 32'h00C64633;
mem['h001A] = 32'h038000EF;
mem['h001B] = 32'h0000006F;
mem['h001C] = 32'h0001A703;
mem['h001D] = 32'h100007B7;
mem['h001E] = 32'h00078793;
mem['h001F] = 32'h00F707B3;
mem['h0020] = 32'h00A70733;
mem['h0021] = 32'h00E1A023;
mem['h0022] = 32'h000016B7;
mem['h0023] = 32'h80068693;
mem['h0024] = 32'h00E6D463;
mem['h0025] = 32'h00100073;
mem['h0026] = 32'h00078513;
mem['h0027] = 32'h00008067;
mem['h0028] = 32'hFD010113;
mem['h0029] = 32'h02400513;
mem['h002A] = 32'h02112623;
mem['h002B] = 32'h02812423;
mem['h002C] = 32'h02912223;
mem['h002D] = 32'h03212023;
mem['h002E] = 32'h01312E23;
mem['h002F] = 32'h01412C23;
mem['h0030] = 32'hFB1FF0EF;
mem['h0031] = 32'h00050413;
mem['h0032] = 32'h00800513;
mem['h0033] = 32'hFA5FF0EF;
mem['h0034] = 32'h00050913;
mem['h0035] = 32'h01C00513;
mem['h0036] = 32'hF99FF0EF;
mem['h0037] = 32'h00050493;
mem['h0038] = 32'h00400513;
mem['h0039] = 32'hF8DFF0EF;
mem['h003A] = 32'h200007B7;
mem['h003B] = 32'h00F52023;
mem['h003C] = 32'h00A4A023;
mem['h003D] = 32'h00400513;
mem['h003E] = 32'hF79FF0EF;
mem['h003F] = 32'h200007B7;
mem['h0040] = 32'h00478793;
mem['h0041] = 32'h00F52023;
mem['h0042] = 32'h00A4A223;
mem['h0043] = 32'h00400513;
mem['h0044] = 32'hF61FF0EF;
mem['h0045] = 32'h200007B7;
mem['h0046] = 32'h00878793;
mem['h0047] = 32'h00F52023;
mem['h0048] = 32'h00A4A423;
mem['h0049] = 32'h00400513;
mem['h004A] = 32'hF49FF0EF;
mem['h004B] = 32'h200007B7;
mem['h004C] = 32'h00C78793;
mem['h004D] = 32'h00F52023;
mem['h004E] = 32'h00A4A623;
mem['h004F] = 32'h00400513;
mem['h0050] = 32'hF31FF0EF;
mem['h0051] = 32'h200007B7;
mem['h0052] = 32'h01078793;
mem['h0053] = 32'h00F52023;
mem['h0054] = 32'h00A4A823;
mem['h0055] = 32'h00400513;
mem['h0056] = 32'hF19FF0EF;
mem['h0057] = 32'h200007B7;
mem['h0058] = 32'h01478793;
mem['h0059] = 32'h00F52023;
mem['h005A] = 32'h00A4AA23;
mem['h005B] = 32'h00400513;
mem['h005C] = 32'hF01FF0EF;
mem['h005D] = 32'h200007B7;
mem['h005E] = 32'h01878793;
mem['h005F] = 32'h00F52023;
mem['h0060] = 32'h00A4AC23;
mem['h0061] = 32'h00992023;
mem['h0062] = 32'h01C00513;
mem['h0063] = 32'hEE5FF0EF;
mem['h0064] = 32'h00050493;
mem['h0065] = 32'h00400513;
mem['h0066] = 32'hED9FF0EF;
mem['h0067] = 32'h200007B7;
mem['h0068] = 32'h01C78793;
mem['h0069] = 32'h00F52023;
mem['h006A] = 32'h00A4A023;
mem['h006B] = 32'h00400513;
mem['h006C] = 32'hEC1FF0EF;
mem['h006D] = 32'h200007B7;
mem['h006E] = 32'h02078793;
mem['h006F] = 32'h00F52023;
mem['h0070] = 32'h00A4A223;
mem['h0071] = 32'h00400513;
mem['h0072] = 32'hEA9FF0EF;
mem['h0073] = 32'h200007B7;
mem['h0074] = 32'h02478793;
mem['h0075] = 32'h00F52023;
mem['h0076] = 32'h00A4A423;
mem['h0077] = 32'h00400513;
mem['h0078] = 32'hE91FF0EF;
mem['h0079] = 32'h200007B7;
mem['h007A] = 32'h02878793;
mem['h007B] = 32'h00F52023;
mem['h007C] = 32'h00A4A623;
mem['h007D] = 32'h00400513;
mem['h007E] = 32'hE79FF0EF;
mem['h007F] = 32'h200007B7;
mem['h0080] = 32'h02C78793;
mem['h0081] = 32'h00F52023;
mem['h0082] = 32'h00A4A823;
mem['h0083] = 32'h00400513;
mem['h0084] = 32'hE61FF0EF;
mem['h0085] = 32'h200007B7;
mem['h0086] = 32'h03078793;
mem['h0087] = 32'h00F52023;
mem['h0088] = 32'h00A4AA23;
mem['h0089] = 32'h00400513;
mem['h008A] = 32'hE49FF0EF;
mem['h008B] = 32'h200007B7;
mem['h008C] = 32'h03478793;
mem['h008D] = 32'h00F52023;
mem['h008E] = 32'h00A4AC23;
mem['h008F] = 32'h00992223;
mem['h0090] = 32'h01242023;
mem['h0091] = 32'h01000513;
mem['h0092] = 32'hE29FF0EF;
mem['h0093] = 32'h00050493;
mem['h0094] = 32'h00400513;
mem['h0095] = 32'hE1DFF0EF;
mem['h0096] = 32'h200007B7;
mem['h0097] = 32'h03878793;
mem['h0098] = 32'h00F52023;
mem['h0099] = 32'h00A4A023;
mem['h009A] = 32'h00400513;
mem['h009B] = 32'hE05FF0EF;
mem['h009C] = 32'h200007B7;
mem['h009D] = 32'h03C78793;
mem['h009E] = 32'h00F52023;
mem['h009F] = 32'h00A4A223;
mem['h00A0] = 32'h00400513;
mem['h00A1] = 32'hDEDFF0EF;
mem['h00A2] = 32'h200007B7;
mem['h00A3] = 32'h04078793;
mem['h00A4] = 32'h00F52023;
mem['h00A5] = 32'h00A4A423;
mem['h00A6] = 32'h00400513;
mem['h00A7] = 32'hDD5FF0EF;
mem['h00A8] = 32'h200007B7;
mem['h00A9] = 32'h04478793;
mem['h00AA] = 32'h00F52023;
mem['h00AB] = 32'h00A4A623;
mem['h00AC] = 32'h00942223;
mem['h00AD] = 32'h00400513;
mem['h00AE] = 32'hDB9FF0EF;
mem['h00AF] = 32'h200007B7;
mem['h00B0] = 32'h04878793;
mem['h00B1] = 32'h00F52023;
mem['h00B2] = 32'h200004B7;
mem['h00B3] = 32'hE0000A37;
mem['h00B4] = 32'h200009B7;
mem['h00B5] = 32'h00A42423;
mem['h00B6] = 32'h04C48493;
mem['h00B7] = 32'hFC0A0A13;
mem['h00B8] = 32'h05C98993;
mem['h00B9] = 32'h00400513;
mem['h00BA] = 32'hD89FF0EF;
mem['h00BB] = 32'h00050913;
mem['h00BC] = 32'h00400513;
mem['h00BD] = 32'hD7DFF0EF;
mem['h00BE] = 32'h00952023;
mem['h00BF] = 32'h014487B3;
mem['h00C0] = 32'h00A92023;
mem['h00C1] = 32'h00F407B3;
mem['h00C2] = 32'h0127A023;
mem['h00C3] = 32'h00448493;
mem['h00C4] = 32'hFD349AE3;
mem['h00C5] = 32'h00400513;
mem['h00C6] = 32'hD59FF0EF;
mem['h00C7] = 32'h00050913;
mem['h00C8] = 32'h00400513;
mem['h00C9] = 32'hD4DFF0EF;
mem['h00CA] = 32'h00952023;
mem['h00CB] = 32'h00A92023;
mem['h00CC] = 32'h01242E23;
mem['h00CD] = 32'h00400513;
mem['h00CE] = 32'hD39FF0EF;
mem['h00CF] = 32'h000F46B7;
mem['h00D0] = 32'h23F68693;
mem['h00D1] = 32'h00842783;
mem['h00D2] = 32'h0007A703;
mem['h00D3] = 32'h00072783;
mem['h00D4] = 32'h2007E793;
mem['h00D5] = 32'h00F72023;
mem['h00D6] = 32'h00842703;
mem['h00D7] = 32'h00842783;
mem['h00D8] = 32'h00072603;
mem['h00D9] = 32'h0007A783;
mem['h00DA] = 32'h0007A703;
mem['h00DB] = 32'h00062783;
mem['h00DC] = 32'h00177713;
mem['h00DD] = 32'h00871713;
mem['h00DE] = 32'hEFF7F793;
mem['h00DF] = 32'h00E7E7B3;
mem['h00E0] = 32'h00F62023;
mem['h00E1] = 32'h00012623;
mem['h00E2] = 32'h00C12783;
mem['h00E3] = 32'h06F6F063;
mem['h00E4] = 32'h00842783;
mem['h00E5] = 32'h0007A703;
mem['h00E6] = 32'h00072783;
mem['h00E7] = 32'hDFF7F793;
mem['h00E8] = 32'h00F72023;
mem['h00E9] = 32'h00842703;
mem['h00EA] = 32'h00842783;
mem['h00EB] = 32'h00072603;
mem['h00EC] = 32'h0007A783;
mem['h00ED] = 32'h0007A703;
mem['h00EE] = 32'h00062783;
mem['h00EF] = 32'h00177713;
mem['h00F0] = 32'h00871713;
mem['h00F1] = 32'hEFF7F793;
mem['h00F2] = 32'h00E7E7B3;
mem['h00F3] = 32'h00F62023;
mem['h00F4] = 32'h00012423;
mem['h00F5] = 32'h00812783;
mem['h00F6] = 32'hF6F6E6E3;
mem['h00F7] = 32'h00812783;
mem['h00F8] = 32'h00178793;
mem['h00F9] = 32'h00F12423;
mem['h00FA] = 32'hFEDFF06F;
mem['h00FB] = 32'h00C12783;
mem['h00FC] = 32'h00178793;
mem['h00FD] = 32'h00F12623;
mem['h00FE] = 32'hF91FF06F;
