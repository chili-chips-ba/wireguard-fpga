-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 6
entity BIN_OP_GT_int17_t_int32_t_0CLK_794ce60a is
port(
 left : in signed(16 downto 0);
 right : in signed(31 downto 0);
 return_output : out unsigned(0 downto 0));
end BIN_OP_GT_int17_t_int32_t_0CLK_794ce60a;
architecture arch of BIN_OP_GT_int17_t_int32_t_0CLK_794ce60a is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- CONST_SR_16[BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912]
signal CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_x : signed(31 downto 0);
signal CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output : signed(31 downto 0);

-- CONST_SR_16[BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1]
signal CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_x : signed(31 downto 0);
signal CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output : signed(31 downto 0);

-- BIN_OP_EQ[BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978]
signal BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_left : unsigned(15 downto 0);
signal BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_right : unsigned(15 downto 0);
signal BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output : unsigned(0 downto 0);

-- rv_MUX[BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9]
signal rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_cond : unsigned(0 downto 0);
signal rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iftrue : unsigned(0 downto 0);
signal rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iffalse : unsigned(0 downto 0);
signal rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output : unsigned(0 downto 0);

-- BIN_OP_GT[BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197]
signal BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_left : unsigned(15 downto 0);
signal BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_right : unsigned(15 downto 0);
signal BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output : unsigned(0 downto 0);

function int32_31_31( x : signed) return unsigned is
--variable x : signed(31 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(31- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912 : 0 clocks latency
CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912 : entity work.CONST_SR_16_int32_t_0CLK_de264c78 port map (
CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_x,
CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output);

-- CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1 : 0 clocks latency
CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1 : entity work.CONST_SR_16_int32_t_0CLK_de264c78 port map (
CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_x,
CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output);

-- BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978 : 0 clocks latency
BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978 : entity work.BIN_OP_EQ_uint16_t_uint16_t_0CLK_de264c78 port map (
BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_left,
BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_right,
BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output);

-- rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9 : 0 clocks latency
rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_cond,
rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iftrue,
rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iffalse,
rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output);

-- BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197 : 0 clocks latency
BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197 : entity work.BIN_OP_GT_uint16_t_uint16_t_0CLK_380ecc95 port map (
BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_left,
BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_right,
BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 left,
 right,
 -- All submodule outputs
 CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output,
 CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output,
 BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output,
 rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output,
 BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_left : signed(16 downto 0);
 variable VAR_right : signed(31 downto 0);
 variable VAR_return_output : unsigned(0 downto 0);
 variable VAR_lsign : unsigned(0 downto 0);
 variable VAR_rsign : unsigned(0 downto 0);
 variable VAR_int32_31_31_BIN_OP_GT_int17_t_int32_t_c_l8_c21_af5d_return_output : unsigned(0 downto 0);
 variable VAR_lsigned : signed(31 downto 0);
 variable VAR_lsigned_BIN_OP_GT_int17_t_int32_t_c_l9_c13_1f23_0 : signed(31 downto 0);
 variable VAR_rsigned : signed(31 downto 0);
 variable VAR_extra_sign_bits : unsigned(15 downto 0);
 variable VAR_extra_sign_bits_BIN_OP_GT_int17_t_int32_t_c_l12_c14_869a_0 : unsigned(15 downto 0);
 variable VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output : signed(31 downto 0);
 variable VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_x : signed(31 downto 0);
 variable VAR_sign_ext_like_zero : unsigned(15 downto 0);
 variable VAR_sign_ext_like_zero_BIN_OP_GT_int17_t_int32_t_c_l13_c14_1408_0 : unsigned(15 downto 0);
 variable VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output : signed(31 downto 0);
 variable VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_x : signed(31 downto 0);
 variable VAR_lunsigned : unsigned(15 downto 0);
 variable VAR_lunsigned_BIN_OP_GT_int17_t_int32_t_c_l16_c14_91e5_0 : unsigned(15 downto 0);
 variable VAR_runsigned : unsigned(15 downto 0);
 variable VAR_runsigned_BIN_OP_GT_int17_t_int32_t_c_l17_c14_d503_0 : unsigned(15 downto 0);
 variable VAR_rv : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output : unsigned(0 downto 0);
 variable VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iftrue : unsigned(0 downto 0);
 variable VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iffalse : unsigned(0 downto 0);
 variable VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output : unsigned(0 downto 0);
 variable VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_left : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_right : unsigned(15 downto 0);
 variable VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_left := left;
     VAR_right := right;

     -- Submodule level 0
     VAR_lsigned_BIN_OP_GT_int17_t_int32_t_c_l9_c13_1f23_0 := resize(VAR_left, 32);
     VAR_lunsigned_BIN_OP_GT_int17_t_int32_t_c_l16_c14_91e5_0 := resize(unsigned(std_logic_vector(VAR_left)),16);
     VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_x := VAR_right;
     VAR_runsigned_BIN_OP_GT_int17_t_int32_t_c_l17_c14_d503_0 := resize(unsigned(std_logic_vector(VAR_right)),16);
     VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_x := VAR_lsigned_BIN_OP_GT_int17_t_int32_t_c_l9_c13_1f23_0;
     VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_left := VAR_lunsigned_BIN_OP_GT_int17_t_int32_t_c_l16_c14_91e5_0;
     VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_right := VAR_runsigned_BIN_OP_GT_int17_t_int32_t_c_l17_c14_d503_0;
     -- CONST_SR_16[BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1] LATENCY=0
     -- Inputs
     CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_x <= VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_x;
     -- Outputs
     VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output := CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output;

     -- CONST_SR_16[BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912] LATENCY=0
     -- Inputs
     CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_x <= VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_x;
     -- Outputs
     VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output := CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output;

     -- int32_31_31[BIN_OP_GT_int17_t_int32_t_c_l8_c21_af5d] LATENCY=0
     VAR_int32_31_31_BIN_OP_GT_int17_t_int32_t_c_l8_c21_af5d_return_output := int32_31_31(
     VAR_right);

     -- BIN_OP_GT[BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197] LATENCY=0
     -- Inputs
     BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_left <= VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_left;
     BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_right <= VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_right;
     -- Outputs
     VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output := BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output;

     -- Submodule level 1
     VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iftrue := VAR_BIN_OP_GT_BIN_OP_GT_int17_t_int32_t_c_l22_c14_d197_return_output;
     VAR_extra_sign_bits_BIN_OP_GT_int17_t_int32_t_c_l12_c14_869a_0 := resize(unsigned(std_logic_vector(VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l12_c32_8912_return_output)),16);
     VAR_sign_ext_like_zero_BIN_OP_GT_int17_t_int32_t_c_l13_c14_1408_0 := resize(unsigned(std_logic_vector(VAR_CONST_SR_16_BIN_OP_GT_int17_t_int32_t_c_l13_c35_11b1_return_output)),16);
     VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iffalse := VAR_int32_31_31_BIN_OP_GT_int17_t_int32_t_c_l8_c21_af5d_return_output;
     VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_left := VAR_extra_sign_bits_BIN_OP_GT_int17_t_int32_t_c_l12_c14_869a_0;
     VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_right := VAR_sign_ext_like_zero_BIN_OP_GT_int17_t_int32_t_c_l13_c14_1408_0;
     -- BIN_OP_EQ[BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978] LATENCY=0
     -- Inputs
     BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_left <= VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_left;
     BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_right <= VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_right;
     -- Outputs
     VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output := BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output;

     -- Submodule level 2
     VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_cond := VAR_BIN_OP_EQ_BIN_OP_GT_int17_t_int32_t_c_l20_c8_7978_return_output;
     -- rv_MUX[BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9] LATENCY=0
     -- Inputs
     rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_cond <= VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_cond;
     rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iftrue <= VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iftrue;
     rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iffalse <= VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_iffalse;
     -- Outputs
     VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output := rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output;

     -- Submodule level 3
     VAR_return_output := VAR_rv_MUX_BIN_OP_GT_int17_t_int32_t_c_l20_c5_27d9_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
