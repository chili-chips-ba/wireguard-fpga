-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 16
entity axis128_keep_count_0CLK_08de2a73 is
port(
 axis : in axis128_t;
 return_output : out unsigned(4 downto 0));
end axis128_keep_count_0CLK_08de2a73;
architecture arch of axis128_keep_count_0CLK_08de2a73 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_d6fa]
signal FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_ae15]
signal FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_e75b]
signal FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_0410]
signal FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_a917]
signal FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_27c7]
signal FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_bf16]
signal FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_26b3]
signal FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_f3f7]
signal FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_8ea0]
signal FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_6f71]
signal FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_9dd0]
signal FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_4697]
signal FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_69ce]
signal FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_03b3]
signal FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_bc25]
signal FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output : unsigned(5 downto 0);


begin

-- SUBMODULE INSTANCES 
-- FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_left,
FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_right,
FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_left,
FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_right,
FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_left,
FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_right,
FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_left,
FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_right,
FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_left,
FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_right,
FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_left,
FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_right,
FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_left,
FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_right,
FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_left,
FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_right,
FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_left,
FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_right,
FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_left,
FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_right,
FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_left,
FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_right,
FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_left,
FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_right,
FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_left,
FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_right,
FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_left,
FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_right,
FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_left,
FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_right,
FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output);

-- FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25 : 0 clocks latency
FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_left,
FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_right,
FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 axis,
 -- All submodule outputs
 FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output,
 FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output,
 FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output,
 FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output,
 FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output,
 FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output,
 FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output,
 FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output,
 FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output,
 FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output,
 FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output,
 FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output,
 FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output,
 FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output,
 FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output,
 FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(4 downto 0);
 variable VAR_axis : axis128_t;
 variable VAR_rv : unsigned(4 downto 0);
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_0_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_1_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_2_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_3_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_4_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_5_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_6_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_7_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_8_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_9_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_10_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_11_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_12_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_13_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_14_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_15_rv_axis_h_l91_c5_33bc : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_4192_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output : unsigned(5 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_left := to_unsigned(0, 5);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_axis := axis;

     -- Submodule level 0
     -- FOR_axis_h_l90_c3_477b_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(7);

     -- FOR_axis_h_l90_c3_477b_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(0);

     -- FOR_axis_h_l90_c3_477b_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(5);

     -- FOR_axis_h_l90_c3_477b_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(14);

     -- FOR_axis_h_l90_c3_477b_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(4);

     -- FOR_axis_h_l90_c3_477b_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(9);

     -- FOR_axis_h_l90_c3_477b_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(11);

     -- FOR_axis_h_l90_c3_477b_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(12);

     -- FOR_axis_h_l90_c3_477b_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(1);

     -- FOR_axis_h_l90_c3_477b_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(2);

     -- FOR_axis_h_l90_c3_477b_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(3);

     -- FOR_axis_h_l90_c3_477b_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(13);

     -- FOR_axis_h_l90_c3_477b_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(8);

     -- FOR_axis_h_l90_c3_477b_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(15);

     -- FOR_axis_h_l90_c3_477b_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(10);

     -- FOR_axis_h_l90_c3_477b_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d[axis_h_l91_c11_4192] LATENCY=0
     VAR_FOR_axis_h_l90_c3_477b_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_4192_return_output := VAR_axis.tkeep(6);

     -- Submodule level 1
     VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_right := VAR_FOR_axis_h_l90_c3_477b_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_right := VAR_FOR_axis_h_l90_c3_477b_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_right := VAR_FOR_axis_h_l90_c3_477b_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_right := VAR_FOR_axis_h_l90_c3_477b_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_right := VAR_FOR_axis_h_l90_c3_477b_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_right := VAR_FOR_axis_h_l90_c3_477b_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_right := VAR_FOR_axis_h_l90_c3_477b_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_right := VAR_FOR_axis_h_l90_c3_477b_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_right := VAR_FOR_axis_h_l90_c3_477b_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_right := VAR_FOR_axis_h_l90_c3_477b_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_right := VAR_FOR_axis_h_l90_c3_477b_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_right := VAR_FOR_axis_h_l90_c3_477b_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_right := VAR_FOR_axis_h_l90_c3_477b_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_right := VAR_FOR_axis_h_l90_c3_477b_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_right := VAR_FOR_axis_h_l90_c3_477b_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_4192_return_output;
     VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_right := VAR_FOR_axis_h_l90_c3_477b_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_4192_return_output;
     -- FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_d6fa] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_left;
     FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output := FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output;

     -- Submodule level 2
     VAR_FOR_axis_h_l90_c3_477b_ITER_0_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_d6fa_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_left := VAR_FOR_axis_h_l90_c3_477b_ITER_0_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_ae15] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_left;
     FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output := FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output;

     -- Submodule level 3
     VAR_FOR_axis_h_l90_c3_477b_ITER_1_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_ae15_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_left := VAR_FOR_axis_h_l90_c3_477b_ITER_1_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_e75b] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_left;
     FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output := FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output;

     -- Submodule level 4
     VAR_FOR_axis_h_l90_c3_477b_ITER_2_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_e75b_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_left := VAR_FOR_axis_h_l90_c3_477b_ITER_2_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_0410] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_left;
     FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output := FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output;

     -- Submodule level 5
     VAR_FOR_axis_h_l90_c3_477b_ITER_3_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_0410_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_left := VAR_FOR_axis_h_l90_c3_477b_ITER_3_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_a917] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_left;
     FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output := FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output;

     -- Submodule level 6
     VAR_FOR_axis_h_l90_c3_477b_ITER_4_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_a917_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_left := VAR_FOR_axis_h_l90_c3_477b_ITER_4_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_27c7] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_left;
     FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output := FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output;

     -- Submodule level 7
     VAR_FOR_axis_h_l90_c3_477b_ITER_5_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_27c7_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_left := VAR_FOR_axis_h_l90_c3_477b_ITER_5_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_bf16] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_left;
     FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output := FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output;

     -- Submodule level 8
     VAR_FOR_axis_h_l90_c3_477b_ITER_6_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_bf16_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_left := VAR_FOR_axis_h_l90_c3_477b_ITER_6_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_26b3] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_left;
     FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output := FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output;

     -- Submodule level 9
     VAR_FOR_axis_h_l90_c3_477b_ITER_7_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_26b3_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_left := VAR_FOR_axis_h_l90_c3_477b_ITER_7_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_f3f7] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_left;
     FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output := FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output;

     -- Submodule level 10
     VAR_FOR_axis_h_l90_c3_477b_ITER_8_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_f3f7_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_left := VAR_FOR_axis_h_l90_c3_477b_ITER_8_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_8ea0] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_left;
     FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output := FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output;

     -- Submodule level 11
     VAR_FOR_axis_h_l90_c3_477b_ITER_9_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_8ea0_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_left := VAR_FOR_axis_h_l90_c3_477b_ITER_9_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_6f71] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_left;
     FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output := FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output;

     -- Submodule level 12
     VAR_FOR_axis_h_l90_c3_477b_ITER_10_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_6f71_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_left := VAR_FOR_axis_h_l90_c3_477b_ITER_10_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_9dd0] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_left;
     FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output := FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output;

     -- Submodule level 13
     VAR_FOR_axis_h_l90_c3_477b_ITER_11_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_9dd0_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_left := VAR_FOR_axis_h_l90_c3_477b_ITER_11_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_4697] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_left;
     FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output := FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output;

     -- Submodule level 14
     VAR_FOR_axis_h_l90_c3_477b_ITER_12_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_4697_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_left := VAR_FOR_axis_h_l90_c3_477b_ITER_12_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_69ce] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_left;
     FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output := FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output;

     -- Submodule level 15
     VAR_FOR_axis_h_l90_c3_477b_ITER_13_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_69ce_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_left := VAR_FOR_axis_h_l90_c3_477b_ITER_13_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_03b3] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_left;
     FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output := FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output;

     -- Submodule level 16
     VAR_FOR_axis_h_l90_c3_477b_ITER_14_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_03b3_return_output, 5);
     VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_left := VAR_FOR_axis_h_l90_c3_477b_ITER_14_rv_axis_h_l91_c5_33bc;
     -- FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_bc25] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_left <= VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_left;
     FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_right <= VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output := FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output;

     -- Submodule level 17
     VAR_FOR_axis_h_l90_c3_477b_ITER_15_rv_axis_h_l91_c5_33bc := resize(VAR_FOR_axis_h_l90_c3_477b_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_bc25_return_output, 5);
     VAR_return_output := VAR_FOR_axis_h_l90_c3_477b_ITER_15_rv_axis_h_l91_c5_33bc;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
