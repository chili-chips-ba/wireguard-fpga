-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 243
entity tb_0CLK_837e73b8 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 global_to_module : in tb_global_to_module_t;
 module_to_global : out tb_module_to_global_t;
 return_output : out axis128_t_stream_t);
end tb_0CLK_837e73b8;
architecture arch of tb_0CLK_837e73b8 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal input_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal ciphertext_in_stream : uint8_t_144 := (others => to_unsigned(0, 8));
signal ciphertext_remaining_in : unsigned(31 downto 0) := to_unsigned(0, 32);
signal cycle_counter : unsigned(31 downto 0) := to_unsigned(0, 32);
signal chacha20poly1305_decrypt_axis_in : axis128_t_stream_t := axis128_t_stream_t_NULL;
signal output_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_size : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_remaining_out : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_expected : char_128 := (others => to_unsigned(0, 8));
signal tag_match_checked : unsigned(0 downto 0) := to_unsigned(0, 1);
signal REG_COMB_input_packet_count : unsigned(31 downto 0);
signal REG_COMB_ciphertext_in_stream : uint8_t_144;
signal REG_COMB_ciphertext_remaining_in : unsigned(31 downto 0);
signal REG_COMB_cycle_counter : unsigned(31 downto 0);
signal REG_COMB_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;
signal REG_COMB_output_packet_count : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_size : unsigned(31 downto 0);
signal REG_COMB_plaintext_remaining_out : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_expected : char_128;
signal REG_COMB_tag_match_checked : unsigned(0 downto 0);

-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l158_c8_2c78]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l159_c1_de5f]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l158_c5_1649]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output : unsigned(31 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l158_c5_1649]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output : uint8_t_144;

-- printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087[chacha20poly1305_decrypt_tb_c_l160_c9_2087]
signal printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087_CLOCK_ENABLE : unsigned(0 downto 0);

-- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l162_c117_5c80]
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_x : unsigned(255 downto 0);
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output : unsigned(255 downto 0);

-- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l162_c148_4c1f]
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_x : unsigned(255 downto 0);
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output : unsigned(255 downto 0);

-- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l162_c179_f337]
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_x : unsigned(255 downto 0);
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output : unsigned(255 downto 0);

-- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l162_c210_b331]
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_x : unsigned(255 downto 0);
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output : unsigned(255 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l162_c241_48be]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_x : unsigned(255 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output : unsigned(255 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l162_c272_22fc]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_x : unsigned(255 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output : unsigned(255 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l162_c302_1732]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_x : unsigned(255 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output : unsigned(255 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l162_c332_0a07]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_x : unsigned(255 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output : unsigned(255 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f[chacha20poly1305_decrypt_tb_c_l162_c64_d73f]
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg3 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg4 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg5 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg6 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg7 : unsigned(31 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l163_c100_db76]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_x : unsigned(95 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output : unsigned(95 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l163_c130_d872]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_x : unsigned(95 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output : unsigned(95 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l163_c160_eb76]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_x : unsigned(95 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output : unsigned(95 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39[chacha20poly1305_decrypt_tb_c_l163_c65_6c39]
signal printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg2 : unsigned(31 downto 0);

-- print_aad[chacha20poly1305_decrypt_tb_c_l164_c9_f355]
signal print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_CLOCK_ENABLE : unsigned(0 downto 0);
signal print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad : uint8_t_32;
signal print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad_len : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l166_c32_54dd]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l167_c35_bdff]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89[chacha20poly1305_decrypt_tb_c_l168_c9_3e89]
signal printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_arg0 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l174_c8_3cb9]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_right : unsigned(0 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l175_c1_53b9]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : unsigned(31 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : unsigned(31 downto 0);

-- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3]
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : axis128_t_stream_t;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : uint8_t_144;

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e]
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);

-- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l186_c56_fbb2]
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_left : unsigned(31 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_right : unsigned(4 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l188_c12_2f43]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l189_c1_747a]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l188_c9_b46a]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output : unsigned(31 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l188_c9_b46a]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output : unsigned(31 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l188_c9_b46a]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output : uint8_t_144;

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l190_c176_7e7d]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l190_c207_b310]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l190_c237_67c4]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l190_c267_bcd3]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98[chacha20poly1305_decrypt_tb_c_l190_c108_ae98]
signal printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg3 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l191_c1_00f0]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l191_c13_99cf]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : unsigned(31 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l191_c13_99cf]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : unsigned(31 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l191_c13_99cf]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : uint8_t_144;

-- printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0[chacha20poly1305_decrypt_tb_c_l192_c17_13c0]
signal printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l194_c17_de27]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output : unsigned(32 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l195_c21_9693]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l196_c1_54a6]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l195_c17_054f]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output : unsigned(31 downto 0);

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l195_c17_054f]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output : uint8_t_144;

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l198_c44_792d]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l199_c47_9bd3]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002[chacha20poly1305_decrypt_tb_c_l200_c21_d002]
signal printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_arg0 : signed(31 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l203_c17_0c24]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l216_c9_8bf0]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l217_c1_17dd]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output : unsigned(0 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : char_128;

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l219_c34_505a]
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_0 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_1 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output : char_array_128_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l220_c30_697f]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68[chacha20poly1305_decrypt_tb_c_l222_c9_cc68]
signal printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_arg0 : unsigned(31 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l228_c8_68e2]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l229_c1_6efc]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : unsigned(31 downto 0);

-- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128]
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : char_128;

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l231_c169_4dfa]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l231_c200_b4b4]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l231_c230_cbe4]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l231_c260_ffc3]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e[chacha20poly1305_decrypt_tb_c_l231_c105_be5e]
signal printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg3 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba]
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l248_c13_209b]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l248_c1_9e99]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf[chacha20poly1305_decrypt_tb_c_l249_c18_8edf]
signal printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_CLOCK_ENABLE : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l252_c1_0b91]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : unsigned(31 downto 0);

-- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364]
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : char_128;

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l253_c16_9d0a]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_right : unsigned(4 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_0e39]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l255_c1_0b96]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : unsigned(31 downto 0);

-- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6]
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : char_128;

-- printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9[chacha20poly1305_decrypt_tb_c_l254_c17_fcd9]
signal printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_CLOCK_ENABLE : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d[chacha20poly1305_decrypt_tb_c_l256_c17_201d]
signal printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_arg0 : signed(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l258_c17_d157]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output : unsigned(32 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l259_c20_173a]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l260_c1_798c]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l259_c17_0f8c]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output : unsigned(31 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l259_c17_0f8c]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l259_c17_0f8c]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output : char_128;

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l262_c43_0b4d]
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_0 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_1 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output : char_array_128_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l264_c42_b292]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3[chacha20poly1305_decrypt_tb_c_l266_c21_57f3]
signal printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_arg0 : signed(31 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l270_c13_ceff]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l276_c5_e2db]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_right : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint8_t_144_uint8_t_144_a26f( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_b938( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;
      base(80) := ref_toks_81;
      base(81) := ref_toks_82;
      base(82) := ref_toks_83;
      base(83) := ref_toks_84;
      base(84) := ref_toks_85;
      base(85) := ref_toks_86;
      base(86) := ref_toks_87;
      base(87) := ref_toks_88;
      base(88) := ref_toks_89;
      base(89) := ref_toks_90;
      base(90) := ref_toks_91;
      base(91) := ref_toks_92;
      base(92) := ref_toks_93;
      base(93) := ref_toks_94;
      base(94) := ref_toks_95;
      base(95) := ref_toks_96;

      return_output := base;
      return return_output; 
end function;

function uint8_array32_be( x : uint8_t_32) return unsigned is

  --variable x : uint8_t_32;
  variable return_output : unsigned(255 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15)&x(16)&x(17)&x(18)&x(19)&x(20)&x(21)&x(22)&x(23)&x(24)&x(25)&x(26)&x(27)&x(28)&x(29)&x(30)&x(31);
return return_output;
end function;

function uint8_array12_be( x : uint8_t_12) return unsigned is

  --variable x : uint8_t_12;
  variable return_output : unsigned(95 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11);
return return_output;
end function;

function CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_16 is
 
  variable base : axis128_t_stream_t; 
  variable return_output : uint8_t_16;
begin
      base.data.tdata(0) := ref_toks_0;
      base.data.tdata(1) := ref_toks_1;
      base.data.tdata(2) := ref_toks_2;
      base.data.tdata(3) := ref_toks_3;
      base.data.tdata(4) := ref_toks_4;
      base.data.tdata(5) := ref_toks_5;
      base.data.tdata(6) := ref_toks_6;
      base.data.tdata(7) := ref_toks_7;
      base.data.tdata(8) := ref_toks_8;
      base.data.tdata(9) := ref_toks_9;
      base.data.tdata(10) := ref_toks_10;
      base.data.tdata(11) := ref_toks_11;
      base.data.tdata(12) := ref_toks_12;
      base.data.tdata(13) := ref_toks_13;
      base.data.tdata(14) := ref_toks_14;
      base.data.tdata(15) := ref_toks_15;

      return_output := base.data.tdata;
      return return_output; 
end function;

function uint8_array16_be( x : uint8_t_16) return unsigned is

  --variable x : uint8_t_16;
  variable return_output : unsigned(127 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15);
return return_output;
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_9fef( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned;
 ref_toks_113 : unsigned;
 ref_toks_114 : unsigned;
 ref_toks_115 : unsigned;
 ref_toks_116 : unsigned;
 ref_toks_117 : unsigned;
 ref_toks_118 : unsigned;
 ref_toks_119 : unsigned;
 ref_toks_120 : unsigned;
 ref_toks_121 : unsigned;
 ref_toks_122 : unsigned;
 ref_toks_123 : unsigned;
 ref_toks_124 : unsigned;
 ref_toks_125 : unsigned;
 ref_toks_126 : unsigned;
 ref_toks_127 : unsigned;
 ref_toks_128 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;
      base(80) := ref_toks_81;
      base(81) := ref_toks_82;
      base(82) := ref_toks_83;
      base(83) := ref_toks_84;
      base(84) := ref_toks_85;
      base(85) := ref_toks_86;
      base(86) := ref_toks_87;
      base(87) := ref_toks_88;
      base(88) := ref_toks_89;
      base(89) := ref_toks_90;
      base(90) := ref_toks_91;
      base(91) := ref_toks_92;
      base(92) := ref_toks_93;
      base(93) := ref_toks_94;
      base(94) := ref_toks_95;
      base(95) := ref_toks_96;
      base(96) := ref_toks_97;
      base(97) := ref_toks_98;
      base(98) := ref_toks_99;
      base(99) := ref_toks_100;
      base(100) := ref_toks_101;
      base(101) := ref_toks_102;
      base(102) := ref_toks_103;
      base(103) := ref_toks_104;
      base(104) := ref_toks_105;
      base(105) := ref_toks_106;
      base(106) := ref_toks_107;
      base(107) := ref_toks_108;
      base(108) := ref_toks_109;
      base(109) := ref_toks_110;
      base(110) := ref_toks_111;
      base(111) := ref_toks_112;
      base(112) := ref_toks_113;
      base(113) := ref_toks_114;
      base(114) := ref_toks_115;
      base(115) := ref_toks_116;
      base(116) := ref_toks_117;
      base(117) := ref_toks_118;
      base(118) := ref_toks_119;
      base(119) := ref_toks_120;
      base(120) := ref_toks_121;
      base(121) := ref_toks_122;
      base(122) := ref_toks_123;
      base(123) := ref_toks_124;
      base(124) := ref_toks_125;
      base(125) := ref_toks_126;
      base(126) := ref_toks_127;
      base(127) := ref_toks_128;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base.data.tkeep(0) := ref_toks_0;
      base.data.tdata(0) := ref_toks_1;
      base.data.tkeep(1) := ref_toks_2;
      base.data.tdata(1) := ref_toks_3;
      base.data.tkeep(2) := ref_toks_4;
      base.data.tdata(2) := ref_toks_5;
      base.data.tkeep(3) := ref_toks_6;
      base.data.tdata(3) := ref_toks_7;
      base.data.tkeep(4) := ref_toks_8;
      base.data.tdata(4) := ref_toks_9;
      base.data.tkeep(5) := ref_toks_10;
      base.data.tdata(5) := ref_toks_11;
      base.data.tkeep(6) := ref_toks_12;
      base.data.tdata(6) := ref_toks_13;
      base.data.tkeep(7) := ref_toks_14;
      base.data.tdata(7) := ref_toks_15;
      base.data.tkeep(8) := ref_toks_16;
      base.data.tdata(8) := ref_toks_17;
      base.data.tkeep(9) := ref_toks_18;
      base.data.tdata(9) := ref_toks_19;
      base.data.tkeep(10) := ref_toks_20;
      base.data.tdata(10) := ref_toks_21;
      base.data.tkeep(11) := ref_toks_22;
      base.data.tdata(11) := ref_toks_23;
      base.data.tkeep(12) := ref_toks_24;
      base.data.tdata(12) := ref_toks_25;
      base.data.tkeep(13) := ref_toks_26;
      base.data.tdata(13) := ref_toks_27;
      base.data.tkeep(14) := ref_toks_28;
      base.data.tdata(14) := ref_toks_29;
      base.data.tkeep(15) := ref_toks_30;
      base.data.tdata(15) := ref_toks_31;
      base.data.tlast := ref_toks_32;
      base.valid := ref_toks_33;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee( ref_toks_0 : axis128_t_stream_t;
 ref_toks_1 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base := ref_toks_0;
      base.valid := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_char_128_char_128_78d0( ref_toks_0 : char_128;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned) return char_128 is
 
  variable base : char_128; 
  variable return_output : char_128;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;
      base(80) := ref_toks_81;
      base(81) := ref_toks_82;
      base(82) := ref_toks_83;
      base(83) := ref_toks_84;
      base(84) := ref_toks_85;
      base(85) := ref_toks_86;
      base(86) := ref_toks_87;
      base(87) := ref_toks_88;
      base(88) := ref_toks_89;
      base(89) := ref_toks_90;
      base(90) := ref_toks_91;
      base(91) := ref_toks_92;
      base(92) := ref_toks_93;
      base(93) := ref_toks_94;
      base(94) := ref_toks_95;
      base(95) := ref_toks_96;
      base(96) := ref_toks_97;
      base(97) := ref_toks_98;
      base(98) := ref_toks_99;
      base(99) := ref_toks_100;
      base(100) := ref_toks_101;
      base(101) := ref_toks_102;
      base(102) := ref_toks_103;
      base(103) := ref_toks_104;
      base(104) := ref_toks_105;
      base(105) := ref_toks_106;
      base(106) := ref_toks_107;
      base(107) := ref_toks_108;
      base(108) := ref_toks_109;
      base(109) := ref_toks_110;
      base(110) := ref_toks_111;
      base(111) := ref_toks_112;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_32_uint8_t_32_1367( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned) return uint8_t_32 is
 
  variable base : uint8_t_32; 
  variable return_output : uint8_t_32;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;
      base(12) := ref_toks_12;
      base(13) := ref_toks_13;
      base(14) := ref_toks_14;
      base(15) := ref_toks_15;
      base(16) := ref_toks_16;
      base(17) := ref_toks_17;
      base(18) := ref_toks_18;
      base(19) := ref_toks_19;
      base(20) := ref_toks_20;
      base(21) := ref_toks_21;
      base(22) := ref_toks_22;
      base(23) := ref_toks_23;
      base(24) := ref_toks_24;
      base(25) := ref_toks_25;
      base(26) := ref_toks_26;
      base(27) := ref_toks_27;
      base(28) := ref_toks_28;
      base(29) := ref_toks_29;
      base(30) := ref_toks_30;
      base(31) := ref_toks_31;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return uint8_t_12 is
 
  variable base : uint8_t_12; 
  variable return_output : uint8_t_12;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78 : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087 : entity work.printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087_CLOCK_ENABLE);

-- CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80 : 0 clocks latency
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80 : entity work.CONST_SR_224_uint256_t_0CLK_de264c78 port map (
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_x,
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output);

-- CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f : 0 clocks latency
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f : entity work.CONST_SR_192_uint256_t_0CLK_de264c78 port map (
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_x,
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output);

-- CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337 : 0 clocks latency
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337 : entity work.CONST_SR_160_uint256_t_0CLK_de264c78 port map (
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_x,
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output);

-- CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331 : 0 clocks latency
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331 : entity work.CONST_SR_128_uint256_t_0CLK_de264c78 port map (
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_x,
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be : entity work.CONST_SR_96_uint256_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc : entity work.CONST_SR_64_uint256_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732 : entity work.CONST_SR_32_uint256_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07 : entity work.CONST_SR_0_uint256_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f : entity work.printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg0,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg1,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg2,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg3,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg4,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg5,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg6,
printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg7);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76 : entity work.CONST_SR_64_uint96_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872 : entity work.CONST_SR_32_uint96_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76 : entity work.CONST_SR_0_uint96_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39 : entity work.printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg0,
printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg1,
printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg2);

-- print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355 : 0 clocks latency
print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355 : entity work.print_aad_0CLK_fa355561 port map (
print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_CLOCK_ENABLE,
print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad,
print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad_len);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89 : entity work.printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_arg0);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9 : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9 : entity work.BIN_OP_GT_uint32_t_uint1_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output);

-- chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : 0 clocks latency
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : entity work.MUX_uint1_t_axis128_t_stream_t_axis128_t_stream_t_0CLK_de264c78 port map (
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

-- BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2 : 0 clocks latency
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2 : entity work.BIN_OP_LTE_uint32_t_uint5_t_0CLK_e595f783 port map (
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_left,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_right,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4 : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3 : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98 : entity work.printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg0,
printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg1,
printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg2,
printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg3);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0 : entity work.printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693 : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693 : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002 : entity work.printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_arg0);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24 : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24 : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0 : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output);

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a : 0 clocks latency
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a : entity work.VAR_REF_RD_char_128_char_2_128_VAR_90b8_0CLK_b45a16e1 port map (
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_1,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_var_dim_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68 : entity work.printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_arg0);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output);

-- output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : 0 clocks latency
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128 : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4 : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3 : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e : entity work.printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg0,
printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg1,
printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg2,
printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg3);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba : entity work.printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf : entity work.printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_CLOCK_ENABLE);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output);

-- output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : 0 clocks latency
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364 : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a : entity work.BIN_OP_GT_uint32_t_uint5_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96 : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output);

-- output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : 0 clocks latency
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6 : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_CLOCK_ENABLE);

-- printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d : entity work.printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output);

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d : 0 clocks latency
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d : entity work.VAR_REF_RD_char_128_char_2_128_VAR_90b8_0CLK_b45a16e1 port map (
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_1,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_var_dim_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3 : entity work.printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_arg0);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334 : 0 clocks latency
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334 : entity work.BIN_OP_MINUS_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_left,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_right,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Registers
 input_packet_count,
 ciphertext_in_stream,
 ciphertext_remaining_in,
 cycle_counter,
 chacha20poly1305_decrypt_axis_in,
 output_packet_count,
 plaintext_out_size,
 plaintext_remaining_out,
 plaintext_out_expected,
 tag_match_checked,
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output,
 CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output,
 CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output,
 CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output,
 CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output,
 chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
 BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output,
 VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output,
 output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output,
 output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output,
 output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output,
 VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output,
 BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_key : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_nonce : uint8_t_12;
 variable VAR_chacha20poly1305_decrypt_aad : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_aad_len : unsigned(7 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out : axis128_t_stream_t;
 variable VAR_key : uint8_t_32;
 variable VAR_nonce : uint8_t_12;
 variable VAR_aad : uint8_t_32;
 variable VAR_aad_len : unsigned(31 downto 0);
 variable VAR_aad_len_chacha20poly1305_decrypt_tb_c_l82_c14_08c0_0 : unsigned(31 downto 0);
 variable VAR_plaintexts : char_2_128;
 variable VAR_plaintext_lens : uint32_t_2;
 variable VAR_input_ciphertext0 : uint8_t_144;
 variable VAR_input_ciphertext1 : uint8_t_144;
 variable VAR_input_ciphertexts : uint8_t_2_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l137_c9_d78f_return_output : uint8_t_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l138_c9_eabc_return_output : uint8_t_144;
 variable VAR_ciphertext_lens : uint32_t_2;
 variable VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l149_c5_0217 : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l166_c9_9c0f : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_PRINT_32_BYTES_uint : unsigned(255 downto 0);
 variable VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg4 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg5 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg6 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg7 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_x : unsigned(255 downto 0);
 variable VAR_PRINT_12_BYTES_uint : unsigned(95 downto 0);
 variable VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l163_c40_3bf0_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_x : unsigned(95 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad : uint8_t_32;
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad_len : unsigned(31 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond : unsigned(0 downto 0);
 variable VAR_i : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond : unsigned(0 downto 0);
 variable VAR_PRINT_16_BYTES_uint : unsigned(127 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l190_c62_4ece_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l190_c45_c0c4_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_x : unsigned(127 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577 : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_144_uint8_t_144_9fef_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l198_c21_6cf3 : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_arg0 : signed(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output : unsigned(31 downto 0);
 variable VAR_ARRAY_SHIFT_DOWN_i : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_16_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_17_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_18_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_19_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_20_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_21_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_22_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_23_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_24_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_25_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_26_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_27_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_28_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_29_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_30_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_31_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_32_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_33_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_34_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_35_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_36_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_37_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_38_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_39_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_40_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_41_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_42_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_43_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_44_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_45_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_46_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_47_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_48_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_49_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_50_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_51_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_52_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_53_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_54_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_55_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_56_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_57_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_58_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_59_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_60_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_61_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_62_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_63_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_64_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_65_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_66_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_67_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_68_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_69_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_70_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_71_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_72_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_73_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_74_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_75_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_76_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_77_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_78_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_79_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_80_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_81_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_82_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_83_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_84_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_85_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_86_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_87_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_88_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_89_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_90_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_91_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_92_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_93_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_94_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_95_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_96_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_97_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_98_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_99_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_100_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_101_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_102_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_103_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_104_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_105_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_106_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_107_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_108_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_109_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_110_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_111_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue : char_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l219_c9_21f1 : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output : char_array_128_t;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_0 : char_128;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_1 : char_128;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l228_c8_2407_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l231_c58_cde3_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l231_c41_722c_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_x : unsigned(127 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_pos : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iffalse : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse : char_128;
 variable VAR_plaintext_out_expected_FALSE_INPUT_MUX_CONST_REF_RD_char_128_char_128_78d0_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : unsigned(31 downto 0);
 variable VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4 : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_arg0 : signed(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue : char_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l262_c18_5b6b : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output : char_array_128_t;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_0 : char_128;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_1 : char_128;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_arg0 : signed(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_0_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_1_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_2_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_3_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_4_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_5_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_6_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_7_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_8_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_9_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_10_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_11_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_12_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_13_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_14_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_15_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_16_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_17_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_18_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_19_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_20_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_21_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_22_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_23_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_24_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_25_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_26_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_27_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_28_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_29_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_30_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_31_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_32_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_33_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_34_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_35_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_36_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_37_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_38_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_39_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_40_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_41_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_42_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_43_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_44_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_45_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_46_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_47_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_48_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_49_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_50_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_51_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_52_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_53_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_54_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_55_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_56_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_57_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_58_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_59_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_60_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_61_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_62_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_63_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_64_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_65_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_66_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_67_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_68_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_69_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_70_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_71_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_72_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_73_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_74_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_75_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_76_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_77_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_78_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_79_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_80_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_81_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_82_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_83_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_84_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_85_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_86_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_87_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_88_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_89_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_90_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_91_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_92_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_93_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_94_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_95_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_96_CONST_REF_RD_char_char_128_112_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_97_CONST_REF_RD_char_char_128_113_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_98_CONST_REF_RD_char_char_128_114_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_99_CONST_REF_RD_char_char_128_115_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_100_CONST_REF_RD_char_char_128_116_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_101_CONST_REF_RD_char_char_128_117_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_102_CONST_REF_RD_char_char_128_118_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_103_CONST_REF_RD_char_char_128_119_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_104_CONST_REF_RD_char_char_128_120_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_105_CONST_REF_RD_char_char_128_121_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_106_CONST_REF_RD_char_char_128_122_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_107_CONST_REF_RD_char_char_128_123_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_108_CONST_REF_RD_char_char_128_124_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_109_CONST_REF_RD_char_char_128_125_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_110_CONST_REF_RD_char_char_128_126_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_111_CONST_REF_RD_char_char_128_127_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output : unsigned(7 downto 0);
 variable VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l276_c5_53b7 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l162_l146_DUPLICATE_b7f0_return_output : uint8_t_32;
 variable VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l147_l163_DUPLICATE_f1d5_return_output : uint8_t_12;
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ecfc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2607_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_11bf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_0aa1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4854_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_8ce5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e021_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ba7d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_bb5e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_3162_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_067d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_f374_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_564f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_10c3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eb68_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_510d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_0911_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_89f4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_d1d3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4cda_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_9d61_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_fe00_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_8cac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eabf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_1186_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e824_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2bd4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_212e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_5494_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_084a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_24c4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_f26a_return_output : unsigned(7 downto 0);
 -- State registers comb logic variables
variable REG_VAR_input_packet_count : unsigned(31 downto 0);
variable REG_VAR_ciphertext_in_stream : uint8_t_144;
variable REG_VAR_ciphertext_remaining_in : unsigned(31 downto 0);
variable REG_VAR_cycle_counter : unsigned(31 downto 0);
variable REG_VAR_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;
variable REG_VAR_output_packet_count : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_size : unsigned(31 downto 0);
variable REG_VAR_plaintext_remaining_out : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_expected : char_128;
variable REG_VAR_tag_match_checked : unsigned(0 downto 0);
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_input_packet_count := input_packet_count;
  REG_VAR_ciphertext_in_stream := ciphertext_in_stream;
  REG_VAR_ciphertext_remaining_in := ciphertext_remaining_in;
  REG_VAR_cycle_counter := cycle_counter;
  REG_VAR_chacha20poly1305_decrypt_axis_in := chacha20poly1305_decrypt_axis_in;
  REG_VAR_output_packet_count := output_packet_count;
  REG_VAR_plaintext_out_size := plaintext_out_size;
  REG_VAR_plaintext_remaining_out := plaintext_remaining_out;
  REG_VAR_plaintext_out_expected := plaintext_out_expected;
  REG_VAR_tag_match_checked := tag_match_checked;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(7, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_right := to_unsigned(0, 1);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_right := to_unsigned(16, 5);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(3, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iffalse := to_unsigned(0, 1);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue := to_unsigned(0, 1);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(6, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_right := to_unsigned(1, 1);
     VAR_chacha20poly1305_decrypt_axis_out_ready := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(13, 32);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_right := to_unsigned(0, 1);
     VAR_chacha20poly1305_decrypt_aad := to_byte_array("Additional authenticated data", 32);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad := to_byte_array("Additional authenticated data", 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(12, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iffalse := to_unsigned(0, 1);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse := to_unsigned(0, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_1 := to_unsigned(71, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_1 := to_unsigned(71, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_1 := to_unsigned(96, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_1 := to_unsigned(96, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iffalse := to_unsigned(0, 1);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(1, 32);
     VAR_aad_len_chacha20poly1305_decrypt_tb_c_l82_c14_08c0_0 := to_unsigned(29, 32);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad_len := VAR_aad_len_chacha20poly1305_decrypt_tb_c_l82_c14_08c0_0;
     VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l149_c5_0217 := resize(VAR_aad_len_chacha20poly1305_decrypt_tb_c_l82_c14_08c0_0, 8);
     VAR_chacha20poly1305_decrypt_aad_len := VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l149_c5_0217;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(11, 32);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(0, 32);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_right := to_unsigned(1, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse := to_unsigned(0, 8);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_0 := to_unsigned(56, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_0 := to_unsigned(56, 32);
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse := to_unsigned(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(15, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(15, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_right := to_unsigned(2, 2);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(15, 32);
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_right := to_unsigned(16, 5);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(5, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_0 := to_unsigned(80, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_0 := to_unsigned(80, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(1, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(1, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_left := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(5, 32);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(2, 32);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_right := to_unsigned(16, 5);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_right := to_unsigned(16, 5);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_right := to_unsigned(2, 2);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right := to_signed(0, 32);
     -- CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l162_l146_DUPLICATE_b7f0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l162_l146_DUPLICATE_b7f0_return_output := CONST_REF_RD_uint8_t_32_uint8_t_32_1367(
     to_unsigned(128, 8),
     to_unsigned(129, 8),
     to_unsigned(130, 8),
     to_unsigned(131, 8),
     to_unsigned(132, 8),
     to_unsigned(133, 8),
     to_unsigned(134, 8),
     to_unsigned(135, 8),
     to_unsigned(136, 8),
     to_unsigned(137, 8),
     to_unsigned(138, 8),
     to_unsigned(139, 8),
     to_unsigned(140, 8),
     to_unsigned(141, 8),
     to_unsigned(142, 8),
     to_unsigned(143, 8),
     to_unsigned(144, 8),
     to_unsigned(145, 8),
     to_unsigned(146, 8),
     to_unsigned(147, 8),
     to_unsigned(148, 8),
     to_unsigned(149, 8),
     to_unsigned(150, 8),
     to_unsigned(151, 8),
     to_unsigned(152, 8),
     to_unsigned(153, 8),
     to_unsigned(154, 8),
     to_unsigned(155, 8),
     to_unsigned(156, 8),
     to_unsigned(157, 8),
     to_unsigned(158, 8),
     to_unsigned(159, 8));

     -- CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l147_l163_DUPLICATE_f1d5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l147_l163_DUPLICATE_f1d5_return_output := CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2(
     to_unsigned(7, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(64, 8),
     to_unsigned(65, 8),
     to_unsigned(66, 8),
     to_unsigned(67, 8),
     to_unsigned(68, 8),
     to_unsigned(69, 8),
     to_unsigned(70, 8),
     to_unsigned(71, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_a26f[chacha20poly1305_decrypt_tb_c_l137_c9_d78f] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l137_c9_d78f_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_a26f(
     (others => to_unsigned(0, 8)),
     to_unsigned(215, 8),
     to_unsigned(30, 8),
     to_unsigned(133, 8),
     to_unsigned(49, 8),
     to_unsigned(110, 8),
     to_unsigned(221, 8),
     to_unsigned(3, 8),
     to_unsigned(242, 8),
     to_unsigned(92, 8),
     to_unsigned(174, 8),
     to_unsigned(198, 8),
     to_unsigned(184, 8),
     to_unsigned(94, 8),
     to_unsigned(232, 8),
     to_unsigned(122, 8),
     to_unsigned(221, 8),
     to_unsigned(225, 8),
     to_unsigned(237, 8),
     to_unsigned(168, 8),
     to_unsigned(104, 8),
     to_unsigned(96, 8),
     to_unsigned(115, 8),
     to_unsigned(11, 8),
     to_unsigned(185, 8),
     to_unsigned(168, 8),
     to_unsigned(235, 8),
     to_unsigned(162, 8),
     to_unsigned(227, 8),
     to_unsigned(117, 8),
     to_unsigned(246, 8),
     to_unsigned(102, 8),
     to_unsigned(196, 8),
     to_unsigned(35, 8),
     to_unsigned(178, 8),
     to_unsigned(235, 8),
     to_unsigned(84, 8),
     to_unsigned(201, 8),
     to_unsigned(250, 8),
     to_unsigned(121, 8),
     to_unsigned(88, 8),
     to_unsigned(152, 8),
     to_unsigned(174, 8),
     to_unsigned(215, 8),
     to_unsigned(124, 8),
     to_unsigned(142, 8),
     to_unsigned(251, 8),
     to_unsigned(38, 8),
     to_unsigned(128, 8),
     to_unsigned(28, 8),
     to_unsigned(119, 8),
     to_unsigned(146, 8),
     to_unsigned(15, 8),
     to_unsigned(219, 8),
     to_unsigned(8, 8),
     to_unsigned(9, 8),
     to_unsigned(110, 8),
     to_unsigned(96, 8),
     to_unsigned(164, 8),
     to_unsigned(133, 8),
     to_unsigned(207, 8),
     to_unsigned(17, 8),
     to_unsigned(184, 8),
     to_unsigned(27, 8),
     to_unsigned(89, 8),
     to_unsigned(93, 8),
     to_unsigned(168, 8),
     to_unsigned(125, 8),
     to_unsigned(106, 8),
     to_unsigned(45, 8),
     to_unsigned(3, 8),
     to_unsigned(201, 8),
     to_unsigned(186, 8),
     to_unsigned(223, 8),
     to_unsigned(92, 8),
     to_unsigned(185, 8),
     to_unsigned(71, 8),
     to_unsigned(116, 8),
     to_unsigned(66, 8),
     to_unsigned(18, 8),
     to_unsigned(63, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_b938[chacha20poly1305_decrypt_tb_c_l138_c9_eabc] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l138_c9_eabc_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_b938(
     (others => to_unsigned(0, 8)),
     to_unsigned(207, 8),
     to_unsigned(18, 8),
     to_unsigned(153, 8),
     to_unsigned(56, 8),
     to_unsigned(109, 8),
     to_unsigned(148, 8),
     to_unsigned(46, 8),
     to_unsigned(223, 8),
     to_unsigned(86, 8),
     to_unsigned(194, 8),
     to_unsigned(230, 8),
     to_unsigned(136, 8),
     to_unsigned(22, 8),
     to_unsigned(245, 8),
     to_unsigned(98, 8),
     to_unsigned(203, 8),
     to_unsigned(225, 8),
     to_unsigned(162, 8),
     to_unsigned(237, 8),
     to_unsigned(76, 8),
     to_unsigned(125, 8),
     to_unsigned(33, 8),
     to_unsigned(38, 8),
     to_unsigned(154, 8),
     to_unsigned(145, 8),
     to_unsigned(170, 8),
     to_unsigned(177, 8),
     to_unsigned(245, 8),
     to_unsigned(58, 8),
     to_unsigned(247, 8),
     to_unsigned(109, 8),
     to_unsigned(193, 8),
     to_unsigned(110, 8),
     to_unsigned(164, 8),
     to_unsigned(226, 8),
     to_unsigned(24, 8),
     to_unsigned(224, 8),
     to_unsigned(235, 8),
     to_unsigned(42, 8),
     to_unsigned(12, 8),
     to_unsigned(203, 8),
     to_unsigned(250, 8),
     to_unsigned(213, 8),
     to_unsigned(96, 8),
     to_unsigned(218, 8),
     to_unsigned(152, 8),
     to_unsigned(26, 8),
     to_unsigned(161, 8),
     to_unsigned(57, 8),
     to_unsigned(77, 8),
     to_unsigned(241, 8),
     to_unsigned(6, 8),
     to_unsigned(215, 8),
     to_unsigned(25, 8),
     to_unsigned(30, 8),
     to_unsigned(111, 8),
     to_unsigned(55, 8),
     to_unsigned(205, 8),
     to_unsigned(247, 8),
     to_unsigned(170, 8),
     to_unsigned(118, 8),
     to_unsigned(205, 8),
     to_unsigned(122, 8),
     to_unsigned(43, 8),
     to_unsigned(152, 8),
     to_unsigned(145, 8),
     to_unsigned(176, 8),
     to_unsigned(58, 8),
     to_unsigned(35, 8),
     to_unsigned(116, 8),
     to_unsigned(207, 8),
     to_unsigned(172, 8),
     to_unsigned(236, 8),
     to_unsigned(106, 8),
     to_unsigned(222, 8),
     to_unsigned(195, 8),
     to_unsigned(78, 8),
     to_unsigned(102, 8),
     to_unsigned(105, 8),
     to_unsigned(120, 8),
     to_unsigned(7, 8),
     to_unsigned(199, 8),
     to_unsigned(227, 8),
     to_unsigned(31, 8),
     to_unsigned(15, 8),
     to_unsigned(235, 8),
     to_unsigned(75, 8),
     to_unsigned(97, 8),
     to_unsigned(234, 8),
     to_unsigned(45, 8),
     to_unsigned(210, 8),
     to_unsigned(164, 8),
     to_unsigned(89, 8),
     to_unsigned(124, 8),
     to_unsigned(174, 8),
     to_unsigned(233, 8));

     -- Submodule level 1
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l138_c9_eabc_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l138_c9_eabc_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l137_c9_d78f_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l137_c9_d78f_return_output;
     VAR_chacha20poly1305_decrypt_nonce := VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l147_l163_DUPLICATE_f1d5_return_output;
     VAR_chacha20poly1305_decrypt_key := VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l162_l146_DUPLICATE_b7f0_return_output;
     -- uint8_array32_be[chacha20poly1305_decrypt_tb_c_l162_c41_b836] LATENCY=0
     VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output := uint8_array32_be(
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l162_l146_DUPLICATE_b7f0_return_output);

     -- uint8_array12_be[chacha20poly1305_decrypt_tb_c_l163_c40_3bf0] LATENCY=0
     VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l163_c40_3bf0_return_output := uint8_array12_be(
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l147_l163_DUPLICATE_f1d5_return_output);

     -- Submodule level 2
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l163_c40_3bf0_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l163_c40_3bf0_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l163_c40_3bf0_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l162_c41_b836_return_output;
     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l162_c302_1732] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l162_c332_0a07] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l163_c100_db76] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output;

     -- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l162_c179_f337] LATENCY=0
     -- Inputs
     CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_x <= VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_x;
     -- Outputs
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output := CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l163_c130_d872] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output;

     -- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l162_c117_5c80] LATENCY=0
     -- Inputs
     CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_x <= VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_x;
     -- Outputs
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output := CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l162_c241_48be] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l163_c160_eb76] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output;

     -- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l162_c148_4c1f] LATENCY=0
     -- Inputs
     CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_x <= VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_x;
     -- Outputs
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output := CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output;

     -- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l162_c210_b331] LATENCY=0
     -- Inputs
     CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_x <= VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_x;
     -- Outputs
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output := CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l162_c272_22fc] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg2 := resize(VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l162_c179_f337_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg3 := resize(VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l162_c210_b331_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg0 := resize(VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l162_c117_5c80_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg2 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l163_c160_eb76_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg4 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l162_c241_48be_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg1 := resize(VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l162_c148_4c1f_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg6 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l162_c302_1732_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg7 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l162_c332_0a07_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg0 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l163_c100_db76_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg5 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l162_c272_22fc_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg1 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l163_c130_d872_return_output, 32);
 -- Reads from global variables
     VAR_chacha20poly1305_decrypt_axis_in_ready := global_to_module.chacha20poly1305_decrypt_axis_in_ready;
     VAR_chacha20poly1305_decrypt_axis_out := global_to_module.chacha20poly1305_decrypt_axis_out;
     -- Submodule level 0
     VAR_return_output := VAR_chacha20poly1305_decrypt_axis_out;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_right := VAR_chacha20poly1305_decrypt_axis_in_ready;
     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eb68 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eb68_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(7);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_067d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_067d_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(5);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_564f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_564f_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(6);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_1186 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_1186_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(12);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_0911 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_0911_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(8);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_9d61 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_9d61_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(10);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_bb5e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_bb5e_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(4);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d[chacha20poly1305_decrypt_tb_c_l228_c8_2407] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l228_c8_2407_return_output := VAR_chacha20poly1305_decrypt_axis_out.valid;

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d[chacha20poly1305_decrypt_tb_c_l231_c58_cde3] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l231_c58_cde3_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4854 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4854_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(2);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_11bf LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_11bf_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(1);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2bd4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2bd4_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(13);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_24c4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_24c4_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(15);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e021 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e021_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(3);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_5494 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_5494_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(14);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d[chacha20poly1305_decrypt_tb_c_l252_c12_fbb3] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tlast;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ecfc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ecfc_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(0);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_8cac LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_8cac_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(11);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_d1d3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_d1d3_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(9);

     -- Submodule level 1
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_24c4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_24c4_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_d1d3_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_d1d3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ecfc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ecfc_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_9d61_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_9d61_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_564f_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_564f_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_left := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l228_c8_2407_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_1186_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_1186_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_bb5e_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_bb5e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_8cac_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_8cac_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_11bf_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_11bf_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_0911_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_0911_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eb68_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eb68_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_067d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_067d_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4854_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4854_return_output, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l252_c12_fbb3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2bd4_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2bd4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e021_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e021_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_5494_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_5494_return_output;
     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l231_c41_722c] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l231_c41_722c_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l231_c58_cde3_return_output);

     -- Submodule level 2
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l231_c41_722c_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l231_c41_722c_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l231_c41_722c_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l231_c41_722c_return_output;
     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l231_c260_ffc3] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l231_c169_4dfa] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l231_c200_b4b4] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l231_c230_cbe4] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l231_c169_4dfa_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l231_c260_ffc3_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l231_c230_cbe4_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l231_c200_b4b4_return_output, 32);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iftrue := VAR_CLOCK_ENABLE;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse := ciphertext_in_stream;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse := ciphertext_remaining_in;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_left := cycle_counter;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_left := input_packet_count;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_var_dim_0 := resize(input_packet_count, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_var_dim_0 := resize(input_packet_count, 1);
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_arg0 := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_arg0 := input_packet_count;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_left := output_packet_count;
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_var_dim_0 := resize(output_packet_count, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_var_dim_0 := resize(output_packet_count, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse := output_packet_count;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse := output_packet_count;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_arg0 := signed(std_logic_vector(resize(output_packet_count, 32)));
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse := plaintext_out_expected;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse := plaintext_out_size;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse := plaintext_remaining_out;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse := tag_match_checked;
     -- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l219_c34_505a] LATENCY=0
     -- Inputs
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_0;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_1 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_ref_toks_1;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_var_dim_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output := VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l216_c9_8bf0] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l158_c8_2c78] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l188_c12_2f43] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l220_c30_697f] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output;

     -- chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee(
     chacha20poly1305_decrypt_axis_in,
     to_unsigned(0, 1));

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l166_c32_54dd] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l228_c8_68e2] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l194_c17_de27] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l258_c17_d157] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l276_c5_e2db] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l167_c35_bdff] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l188_c12_2f43_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l228_c8_68e2_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l158_c8_2c78_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l216_c9_8bf0_return_output;
     VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l194_c17_de27_return_output, 32);
     VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l258_c17_d157_return_output, 32);
     VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l276_c5_53b7 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l276_c5_e2db_return_output, 32);
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l219_c9_21f1 := VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l219_c34_505a_return_output.data;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l167_c35_bdff_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l220_c30_697f_return_output;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l166_c9_9c0f := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l166_c32_54dd_return_output.data;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse := VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l166_c9_9c0f;
     REG_VAR_cycle_counter := VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l276_c5_53b7;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_left := VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_var_dim_0 := resize(VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_var_dim_0 := resize(VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577, 1);
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue := VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_arg0 := signed(std_logic_vector(resize(VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l194_c17_d577, 32)));
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_left := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4;
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_arg0 := signed(std_logic_vector(resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l258_c17_b7c4, 32)));
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l219_c9_21f1;
     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l264_c42_b292] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l199_c47_9bd3] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l158_c5_1649] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l159_c1_de5f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l217_c1_17dd] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l259_c20_173a] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l158_c5_1649] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l198_c44_792d] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output;

     -- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l262_c43_0b4d] LATENCY=0
     -- Inputs
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_0;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_1 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_ref_toks_1;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_var_dim_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output := VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l216_c5_92ea] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l195_c21_9693] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l229_c1_6efc] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;

     -- Submodule level 2
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l195_c21_9693_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l259_c20_173a_return_output;
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l159_c1_de5f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_17dd_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l229_c1_6efc_return_output;
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l262_c18_5b6b := VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l262_c43_0b4d_return_output.data;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l199_c47_9bd3_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l264_c42_b292_return_output;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l198_c21_6cf3 := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l198_c44_792d_return_output.data;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output, 33)));
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_left := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_right := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output, 33)));
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     REG_VAR_tag_match_checked := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l198_c21_6cf3;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l262_c18_5b6b;
     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l248_c13_209b] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_59_CONST_REF_RD_char_char_128_75_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_59_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(75);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_106_CONST_REF_RD_char_char_128_122_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_106_CONST_REF_RD_char_char_128_122_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(122);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(143);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_79_CONST_REF_RD_char_char_128_95_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_79_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(95);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_76_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_76_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(92);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_48_CONST_REF_RD_char_char_128_64_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_48_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(64);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_17_CONST_REF_RD_char_char_128_33_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_17_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(33);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_44_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_44_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(60);

     -- printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087[chacha20poly1305_decrypt_tb_c_l160_c9_2087] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l160_c9_2087_chacha20poly1305_decrypt_tb_c_l160_c9_2087_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_28_CONST_REF_RD_char_char_128_44_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_28_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(44);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_83_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_83_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(99);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_58_CONST_REF_RD_char_char_128_74_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_58_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(74);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(2);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_42_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_42_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(58);

     -- CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_f374 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_f374_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(5);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_64_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_64_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(80);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l203_c17_0c24] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_6_CONST_REF_RD_char_char_128_22_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_6_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(22);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_61_CONST_REF_RD_char_char_128_77_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_61_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(77);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_2_CONST_REF_RD_char_char_128_18_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_2_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(18);

     -- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334 LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_left <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_left;
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_right <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output := BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(11);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(30);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_47_CONST_REF_RD_char_char_128_63_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_47_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(63);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_110_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_110_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(126);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_96_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_96_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(112);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(22);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_103_CONST_REF_RD_char_char_128_119_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_103_CONST_REF_RD_char_char_128_119_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(119);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_16_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_16_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(32);

     -- CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_510d LATENCY=0
     VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_510d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(7);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_37_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_37_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(53);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(139);

     -- CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eabf LATENCY=0
     VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eabf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(11);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_10_CONST_REF_RD_char_char_128_26_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_10_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(26);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(0);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_109_CONST_REF_RD_char_char_128_125_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_109_CONST_REF_RD_char_char_128_125_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(125);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(7);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(136);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_70_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_70_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(86);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_31_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_31_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(47);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_85_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_85_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(101);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_88_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_88_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(104);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l174_c8_3cb9] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_109_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_109_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(125);

     -- printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f[chacha20poly1305_decrypt_tb_c_l162_c64_d73f] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg3;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg4 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg4;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg5 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg5;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg6 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg6;
     printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg7 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_chacha20poly1305_decrypt_tb_c_l162_c64_d73f_arg7;
     -- Outputs

     -- CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_fe00 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_fe00_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(10);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(134);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_39_CONST_REF_RD_char_char_128_55_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_39_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(55);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_9_CONST_REF_RD_char_char_128_25_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_9_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(25);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_0_CONST_REF_RD_char_char_128_16_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_0_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(16);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_32_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_32_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(48);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_7_CONST_REF_RD_char_char_128_23_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_7_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(23);

     -- CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e824 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e824_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(12);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(142);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_44_CONST_REF_RD_char_char_128_60_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_44_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(60);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_97_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_97_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(113);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_80_CONST_REF_RD_char_char_128_96_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_80_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(96);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(9);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_84_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_84_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(100);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_66_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_66_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(82);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_30_CONST_REF_RD_char_char_128_46_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_30_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(46);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_22_CONST_REF_RD_char_char_128_38_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_22_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(38);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_27_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_27_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(43);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(133);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_52_CONST_REF_RD_char_char_128_68_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_52_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(68);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_56_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_56_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(72);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_41_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_41_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(57);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_92_CONST_REF_RD_char_char_128_108_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_92_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(108);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_62_CONST_REF_RD_char_char_128_78_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_62_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(78);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_29_CONST_REF_RD_char_char_128_45_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_29_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(45);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_24_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_24_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(40);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_93_CONST_REF_RD_char_char_128_109_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_93_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(109);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_97_CONST_REF_RD_char_char_128_113_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_97_CONST_REF_RD_char_char_128_113_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(113);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_89_CONST_REF_RD_char_char_128_105_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_89_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(105);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_103_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_103_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(119);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(20);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_53_CONST_REF_RD_char_char_128_69_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_53_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(69);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_76_CONST_REF_RD_char_char_128_92_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_76_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(92);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_21_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_21_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(37);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(31);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(25);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_25_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_25_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(41);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_89_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_89_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(105);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_21_CONST_REF_RD_char_char_128_37_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_21_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(37);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_99_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_99_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(115);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_34_CONST_REF_RD_char_char_128_50_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_34_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(50);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_19_CONST_REF_RD_char_char_128_35_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_19_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(35);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_50_CONST_REF_RD_char_char_128_66_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_50_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(66);

     -- CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_3162 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_3162_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(4);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_65_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_65_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(81);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_31_CONST_REF_RD_char_char_128_47_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_31_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(47);

     -- CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ba7d LATENCY=0
     VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ba7d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(3);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_87_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_87_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(103);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_61_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_61_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(77);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_92_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_92_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(108);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(135);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(18);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_93_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_93_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(109);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_81_CONST_REF_RD_char_char_128_97_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_81_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(97);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_46_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_46_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(62);

     -- CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_0aa1 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_0aa1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(1);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_63_CONST_REF_RD_char_char_128_79_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_63_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(79);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(14);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_67_CONST_REF_RD_char_char_128_83_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_67_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(83);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_81_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_81_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(97);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(28);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_111_CONST_REF_RD_char_char_128_127_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_111_CONST_REF_RD_char_char_128_127_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(127);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_108_CONST_REF_RD_char_char_128_124_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_108_CONST_REF_RD_char_char_128_124_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(124);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l259_c17_0f8c] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(130);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_57_CONST_REF_RD_char_char_128_73_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_57_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(73);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_75_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_75_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(91);

     -- print_aad[chacha20poly1305_decrypt_tb_c_l164_c9_f355] LATENCY=0
     -- Clock enable
     print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_CLOCK_ENABLE <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_CLOCK_ENABLE;
     -- Inputs
     print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad;
     print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad_len <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l164_c9_f355_aad_len;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68[chacha20poly1305_decrypt_tb_c_l222_c9_cc68] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_chacha20poly1305_decrypt_tb_c_l222_c9_cc68_arg0;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_48_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_48_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(64);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_108_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_108_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(124);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_79_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_79_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(95);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_5_CONST_REF_RD_char_char_128_21_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_5_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(21);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_77_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_77_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(93);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_45_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_45_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(61);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(137);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_73_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_73_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(89);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(8);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_54_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_54_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(70);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_73_CONST_REF_RD_char_char_128_89_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_73_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(89);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_57_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_57_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(73);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_72_CONST_REF_RD_char_char_128_88_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_72_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(88);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_65_CONST_REF_RD_char_char_128_81_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_65_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(81);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_90_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_90_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(106);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_86_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_86_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(102);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_12_CONST_REF_RD_char_char_128_28_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_12_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(28);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_42_CONST_REF_RD_char_char_128_58_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_42_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(58);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_75_CONST_REF_RD_char_char_128_91_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_75_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(91);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_47_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_47_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(63);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_29_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_29_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(45);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_85_CONST_REF_RD_char_char_128_101_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_85_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(101);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l195_c17_054f] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_28_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_28_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(44);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_70_CONST_REF_RD_char_char_128_86_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_70_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(86);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_96_CONST_REF_RD_char_char_128_112_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_96_CONST_REF_RD_char_char_128_112_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(112);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_46_CONST_REF_RD_char_char_128_62_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_46_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(62);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_33_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_33_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(49);

     -- printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89[chacha20poly1305_decrypt_tb_c_l168_c9_3e89] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_chacha20poly1305_decrypt_tb_c_l168_c9_3e89_arg0;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_40_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_40_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(56);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(17);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_110_CONST_REF_RD_char_char_128_126_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_110_CONST_REF_RD_char_char_128_126_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(126);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_51_CONST_REF_RD_char_char_128_67_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_51_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(67);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(23);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_91_CONST_REF_RD_char_char_128_107_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_91_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(107);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_39_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_39_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(55);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_78_CONST_REF_RD_char_char_128_94_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_78_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(94);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_94_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_94_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(110);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(21);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_71_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_71_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(87);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_23_CONST_REF_RD_char_char_128_39_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_23_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(39);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_82_CONST_REF_RD_char_char_128_98_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_82_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(98);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_101_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_101_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(117);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(10);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(3);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_100_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_100_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(116);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(13);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_36_CONST_REF_RD_char_char_128_52_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_36_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(52);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_64_CONST_REF_RD_char_char_128_80_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_64_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(80);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_20_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_20_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(36);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_68_CONST_REF_RD_char_char_128_84_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_68_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(84);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_24_CONST_REF_RD_char_char_128_40_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_24_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(40);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(140);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(1);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_95_CONST_REF_RD_char_char_128_111_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_95_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(111);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_86_CONST_REF_RD_char_char_128_102_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_86_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(102);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_104_CONST_REF_RD_char_char_128_120_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_104_CONST_REF_RD_char_char_128_120_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(120);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(19);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_3_CONST_REF_RD_char_char_128_19_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_3_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(19);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_80_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_80_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(96);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_101_CONST_REF_RD_char_char_128_117_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_101_CONST_REF_RD_char_char_128_117_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(117);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_98_CONST_REF_RD_char_char_128_114_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_98_CONST_REF_RD_char_char_128_114_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(114);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(128);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_11_CONST_REF_RD_char_char_128_27_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_11_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(27);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_26_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_26_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(42);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_18_CONST_REF_RD_char_char_128_34_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_18_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(34);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(132);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_16_CONST_REF_RD_char_char_128_32_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_16_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(32);

     -- CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4cda LATENCY=0
     VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4cda_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(9);

     -- CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_212e LATENCY=0
     VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_212e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(13);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_111_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_111_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(127);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_54_CONST_REF_RD_char_char_128_70_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_54_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(70);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_23_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_23_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(39);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_84_CONST_REF_RD_char_char_128_100_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_84_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(100);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_60_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_60_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(76);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_26_CONST_REF_RD_char_char_128_42_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_26_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(42);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_38_CONST_REF_RD_char_char_128_54_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_38_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(54);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_99_CONST_REF_RD_char_char_128_115_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_99_CONST_REF_RD_char_char_128_115_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(115);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l195_c17_054f] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_37_CONST_REF_RD_char_char_128_53_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_37_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(53);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_105_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_105_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(121);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_18_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_18_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(34);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_67_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_67_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(83);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_102_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_102_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(118);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_74_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_74_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(90);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_50_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_50_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(66);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_68_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_68_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(84);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_83_CONST_REF_RD_char_char_128_99_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_83_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(99);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_4_CONST_REF_RD_char_char_128_20_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_4_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(20);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_69_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_69_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(85);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_33_CONST_REF_RD_char_char_128_49_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_33_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(49);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_30_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_30_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(46);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(26);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_87_CONST_REF_RD_char_char_128_103_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_87_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(103);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_22_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_22_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(38);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(27);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_1_CONST_REF_RD_char_char_128_17_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_1_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(17);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_27_CONST_REF_RD_char_char_128_43_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_27_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(43);

     -- CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_10c3 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_10c3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(6);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_107_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_107_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(123);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_82_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_82_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(98);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_58_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_58_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(74);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_38_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_38_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(54);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_51_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_51_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(67);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_63_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_63_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(79);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_8_CONST_REF_RD_char_char_128_24_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_8_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(24);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_100_CONST_REF_RD_char_char_128_116_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_100_CONST_REF_RD_char_char_128_116_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(116);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_55_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_55_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(71);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(141);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_72_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_72_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(88);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_78_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_78_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(94);

     -- printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e[chacha20poly1305_decrypt_tb_c_l231_c105_be5e] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_chacha20poly1305_decrypt_tb_c_l231_c105_be5e_arg3;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_43_CONST_REF_RD_char_char_128_59_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_43_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(59);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_19_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_19_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(35);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_13_CONST_REF_RD_char_char_128_29_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_13_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(29);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2607 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2607_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(0);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_35_CONST_REF_RD_char_char_128_51_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_35_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(51);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_59_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_59_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(75);

     -- CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_f26a LATENCY=0
     VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_f26a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(15);

     -- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l186_c56_fbb2] LATENCY=0
     -- Inputs
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_left <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_left;
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_right <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_right;
     -- Outputs
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output := BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_49_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_49_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(65);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_90_CONST_REF_RD_char_char_128_106_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_90_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(106);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_35_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_35_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(51);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_95_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_95_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(111);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_52_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_52_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(68);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_53_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_53_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(69);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(12);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(129);

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l259_c17_0f8c] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_107_CONST_REF_RD_char_char_128_123_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_107_CONST_REF_RD_char_char_128_123_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(123);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_17_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_17_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(33);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(4);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(5);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_43_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_43_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(59);

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l259_c17_0f8c] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_66_CONST_REF_RD_char_char_128_82_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_66_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(82);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_88_CONST_REF_RD_char_char_128_104_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_88_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(104);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_20_CONST_REF_RD_char_char_128_36_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_20_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(36);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_62_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_62_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(78);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_41_CONST_REF_RD_char_char_128_57_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_41_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(57);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_14_CONST_REF_RD_char_char_128_30_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_14_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(30);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(24);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_55_CONST_REF_RD_char_char_128_71_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_55_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(71);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(15);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_49_CONST_REF_RD_char_char_128_65_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_49_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(65);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_77_CONST_REF_RD_char_char_128_93_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_77_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(93);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_45_CONST_REF_RD_char_char_128_61_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_45_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(61);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_69_CONST_REF_RD_char_char_128_85_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_69_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(85);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_36_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_36_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(52);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l270_c13_ceff] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(131);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_15_CONST_REF_RD_char_char_128_31_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_15_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(31);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_60_CONST_REF_RD_char_char_128_76_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_60_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(76);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_74_CONST_REF_RD_char_char_128_90_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_74_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(90);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_102_CONST_REF_RD_char_char_128_118_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_102_CONST_REF_RD_char_char_128_118_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(118);

     -- CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_084a LATENCY=0
     VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_084a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(14);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(16);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_104_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_104_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(120);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_94_CONST_REF_RD_char_char_128_110_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_94_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(110);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_40_CONST_REF_RD_char_char_128_56_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_40_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(56);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_25_CONST_REF_RD_char_char_128_41_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_25_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(41);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(138);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_98_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_98_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(114);

     -- CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_8ce5 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_8ce5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(2);

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l252_c1_0b91] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_34_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_34_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(50);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l236_c16_29a5] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_56_CONST_REF_RD_char_char_128_72_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_56_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(72);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l181_c16_ff6d] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_left;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d[chacha20poly1305_decrypt_tb_c_l183_c66_56c5] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(6);

     -- printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39[chacha20poly1305_decrypt_tb_c_l163_c65_6c39] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_chacha20poly1305_decrypt_tb_c_l163_c65_6c39_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_71_CONST_REF_RD_char_char_128_87_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_71_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(87);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_106_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_106_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(122);

     -- CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_89f4 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_89f4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(8);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_105_CONST_REF_RD_char_char_128_121_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_105_CONST_REF_RD_char_char_128_121_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(121);

     -- FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_32_CONST_REF_RD_char_char_128_48_d41d[chacha20poly1305_decrypt_tb_c_l271_c164_08b3] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_32_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output(48);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_91_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_91_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(107);

     -- FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d[chacha20poly1305_decrypt_tb_c_l204_c173_59d9] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output(29);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l253_c16_9d0a] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l248_c13_209b_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l174_c8_3cb9_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l253_c16_9d0a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l203_c17_0c24_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l270_c13_ceff_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l240_DUPLICATE_e334_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2607_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_2607_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_fe00_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_fe00_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eabf_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_eabf_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e824_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_e824_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_212e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_212e_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_084a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_084a_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_f26a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_f26a_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_0aa1_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_0aa1_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_8ce5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_8ce5_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ba7d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_ba7d_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_3162_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_3162_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_f374_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_f374_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_10c3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_10c3_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_510d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_510d_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_89f4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l242_l238_DUPLICATE_89f4_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right := VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4cda_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 := resize(VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l238_l242_DUPLICATE_4cda_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l181_c16_ff6d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l183_c66_56c5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l236_c16_29a5_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l252_c1_0b91_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l195_c17_054f_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l259_c17_0f8c_return_output;
     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6] LATENCY=0
     -- Inputs
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse;
     -- Outputs
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output := output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;

     -- plaintext_out_expected_FALSE_INPUT_MUX_CONST_REF_RD_char_128_char_128_78d0[chacha20poly1305_decrypt_tb_c_l252_c9_0364] LATENCY=0
     VAR_plaintext_out_expected_FALSE_INPUT_MUX_CONST_REF_RD_char_128_char_128_78d0_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output := CONST_REF_RD_char_128_char_128_78d0(
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l216_c5_92ea_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_0_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_1_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_2_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_3_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_4_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_5_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_6_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_7_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_8_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_9_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_10_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_11_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_12_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_13_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_14_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_15_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_16_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_17_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_18_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_19_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_20_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_21_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_22_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_23_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_24_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_25_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_26_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_27_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_28_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_29_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_30_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_31_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_32_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_33_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_34_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_35_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_36_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_37_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_38_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_39_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_40_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_41_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_42_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_43_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_44_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_45_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_46_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_47_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_48_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_49_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_50_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_51_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_52_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_53_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_54_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_55_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_56_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_57_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_58_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_59_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_60_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_61_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_62_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_63_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_64_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_65_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_66_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_67_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_68_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_69_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_70_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_71_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_72_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_73_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_74_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_75_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_76_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_77_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_78_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_79_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_80_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_81_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_82_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_83_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_84_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_85_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_86_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_87_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_88_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_89_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_90_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_91_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_92_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_93_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_94_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_95_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_96_CONST_REF_RD_char_char_128_112_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_97_CONST_REF_RD_char_char_128_113_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_98_CONST_REF_RD_char_char_128_114_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_99_CONST_REF_RD_char_char_128_115_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_100_CONST_REF_RD_char_char_128_116_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_101_CONST_REF_RD_char_char_128_117_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_102_CONST_REF_RD_char_char_128_118_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_103_CONST_REF_RD_char_char_128_119_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_104_CONST_REF_RD_char_char_128_120_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_105_CONST_REF_RD_char_char_128_121_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_106_CONST_REF_RD_char_char_128_122_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_107_CONST_REF_RD_char_char_128_123_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_108_CONST_REF_RD_char_char_128_124_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_109_CONST_REF_RD_char_char_128_125_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_110_CONST_REF_RD_char_char_128_126_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l271_c42_fb09_ITER_111_CONST_REF_RD_char_char_128_127_d41d_chacha20poly1305_decrypt_tb_c_l271_c164_08b3_return_output);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l253_c1_0e39] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l191_c13_99cf] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;

     -- ciphertext_in_stream_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_144_uint8_t_144_9fef[chacha20poly1305_decrypt_tb_c_l191_c13_99cf] LATENCY=0
     VAR_ciphertext_in_stream_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_144_uint8_t_144_9fef_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_9fef(
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l158_c5_1649_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_0_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_1_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_2_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_3_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_4_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_5_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_6_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_7_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_8_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_9_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_10_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_11_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_12_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_13_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_14_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_15_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_16_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_17_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_18_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_19_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_20_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_21_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_22_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_23_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_24_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_25_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_26_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_27_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_28_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_29_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_30_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_31_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_32_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_33_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_34_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_35_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_36_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_37_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_38_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_39_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_40_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_41_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_42_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_43_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_44_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_45_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_46_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_47_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_48_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_49_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_50_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_51_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_52_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_53_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_54_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_55_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_56_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_57_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_58_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_59_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_60_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_61_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_62_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_63_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_64_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_65_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_66_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_67_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_68_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_69_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_70_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_71_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_72_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_73_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_74_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_75_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_76_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_77_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_78_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_79_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_80_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_81_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_82_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_83_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_84_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_85_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_86_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_87_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_88_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_89_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_90_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_91_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_92_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_93_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_94_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_95_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_96_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_97_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_98_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_99_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_100_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_101_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_102_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_103_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_104_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_105_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_106_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_107_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_108_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_109_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_110_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_111_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l204_c46_a095_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l204_c173_59d9_return_output);

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l255_c1_0b96] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l253_c13_40a6] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l175_c1_53b9] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l191_c13_99cf] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l248_c1_9e99] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l181_c13_325e] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output := FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l240_c47_eac1] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l237_c1_d6e7] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l238_c20_fc9c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_left;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;

     -- Submodule level 4
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_0b96_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l238_c20_fc9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l240_c47_eac1_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l237_c1_d6e7_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l175_c1_53b9_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l248_c1_9e99_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l253_c1_0e39_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse := VAR_ciphertext_in_stream_FALSE_INPUT_MUX_CONST_REF_RD_uint8_t_144_uint8_t_144_9fef_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse := VAR_plaintext_out_expected_FALSE_INPUT_MUX_CONST_REF_RD_char_128_char_128_78d0_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l253_c13_40a6_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l240_c30_df6a_0;
     -- chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c(
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l186_c56_fbb2_return_output,
     to_unsigned(1, 1));

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l260_c1_798c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9[chacha20poly1305_decrypt_tb_c_l254_c17_fcd9] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_chacha20poly1305_decrypt_tb_c_l254_c17_fcd9_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d[chacha20poly1305_decrypt_tb_c_l256_c17_201d] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_201d_chacha20poly1305_decrypt_tb_c_l256_c17_201d_arg0;
     -- Outputs

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l188_c9_b46a] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed[chacha20poly1305_decrypt_tb_c_l190_c62_4ece] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l190_c62_4ece_return_output := CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed(
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l177_c9_01c8_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l181_c13_325e_return_output);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf[chacha20poly1305_decrypt_tb_c_l249_c18_8edf] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_chacha20poly1305_decrypt_tb_c_l249_c18_8edf_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l188_c9_b46a] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l239_c1_741c] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output := FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l191_c13_99cf] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;

     -- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l252_c9_0364] LATENCY=0
     -- Inputs
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_cond;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iftrue;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_iffalse;
     -- Outputs
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output := output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l189_c1_747a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output;

     -- Submodule level 5
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l239_c1_741c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l189_c1_747a_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l260_c1_798c_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue := VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l191_c13_99cf_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l252_c9_0364_return_output;
     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;

     -- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3] LATENCY=0
     -- Inputs
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse;
     -- Outputs
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output := chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;

     -- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128] LATENCY=0
     -- Inputs
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse;
     -- Outputs
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output := output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l188_c9_b46a] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3[chacha20poly1305_decrypt_tb_c_l266_c21_57f3] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_chacha20poly1305_decrypt_tb_c_l266_c21_57f3_arg0;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l191_c1_00f0] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l190_c45_c0c4] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l190_c45_c0c4_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l190_c62_4ece_return_output);

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l228_c5_6128] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba[chacha20poly1305_decrypt_tb_c_l241_c21_feba] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l234_c9_8fd3_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l241_c21_feba_chacha20poly1305_decrypt_tb_c_l241_c21_feba_arg2;
     -- Outputs

     -- Submodule level 6
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l191_c1_00f0_return_output;
     REG_VAR_chacha20poly1305_decrypt_axis_in := VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l188_c9_b46a_return_output;
     REG_VAR_ciphertext_remaining_in := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;
     REG_VAR_input_packet_count := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;
     REG_VAR_output_packet_count := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;
     REG_VAR_plaintext_out_expected := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;
     REG_VAR_plaintext_out_size := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;
     REG_VAR_plaintext_remaining_out := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l228_c5_6128_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l190_c45_c0c4_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l190_c45_c0c4_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l190_c45_c0c4_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l190_c45_c0c4_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l196_c1_54a6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l190_c237_67c4] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0[chacha20poly1305_decrypt_tb_c_l192_c17_13c0] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_chacha20poly1305_decrypt_tb_c_l192_c17_13c0_arg0;
     -- Outputs

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l174_c5_8dd3] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l190_c267_bcd3] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l190_c176_7e7d] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l190_c207_b310] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output;

     -- Submodule level 7
     VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l190_c267_bcd3_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l190_c237_67c4_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l190_c207_b310_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l190_c176_7e7d_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l196_c1_54a6_return_output;
     REG_VAR_ciphertext_in_stream := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l174_c5_8dd3_return_output;
     -- printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002[chacha20poly1305_decrypt_tb_c_l200_c21_d002] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l200_c21_d002_chacha20poly1305_decrypt_tb_c_l200_c21_d002_arg0;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98[chacha20poly1305_decrypt_tb_c_l190_c108_ae98] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_chacha20poly1305_decrypt_tb_c_l190_c108_ae98_arg3;
     -- Outputs

     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_input_packet_count <= REG_VAR_input_packet_count;
REG_COMB_ciphertext_in_stream <= REG_VAR_ciphertext_in_stream;
REG_COMB_ciphertext_remaining_in <= REG_VAR_ciphertext_remaining_in;
REG_COMB_cycle_counter <= REG_VAR_cycle_counter;
REG_COMB_chacha20poly1305_decrypt_axis_in <= REG_VAR_chacha20poly1305_decrypt_axis_in;
REG_COMB_output_packet_count <= REG_VAR_output_packet_count;
REG_COMB_plaintext_out_size <= REG_VAR_plaintext_out_size;
REG_COMB_plaintext_remaining_out <= REG_VAR_plaintext_remaining_out;
REG_COMB_plaintext_out_expected <= REG_VAR_plaintext_out_expected;
REG_COMB_tag_match_checked <= REG_VAR_tag_match_checked;
-- Global wires driven various places in pipeline
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_key <= VAR_chacha20poly1305_decrypt_key;
else
  module_to_global.chacha20poly1305_decrypt_key <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_nonce <= VAR_chacha20poly1305_decrypt_nonce;
else
  module_to_global.chacha20poly1305_decrypt_nonce <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad <= VAR_chacha20poly1305_decrypt_aad;
else
  module_to_global.chacha20poly1305_decrypt_aad <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad_len <= VAR_chacha20poly1305_decrypt_aad_len;
else
  module_to_global.chacha20poly1305_decrypt_aad_len <= to_unsigned(0, 8);
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= VAR_chacha20poly1305_decrypt_axis_out_ready;
else
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= to_unsigned(0, 1);
end if;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     input_packet_count <= REG_COMB_input_packet_count;
     ciphertext_in_stream <= REG_COMB_ciphertext_in_stream;
     ciphertext_remaining_in <= REG_COMB_ciphertext_remaining_in;
     cycle_counter <= REG_COMB_cycle_counter;
     chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in;
     output_packet_count <= REG_COMB_output_packet_count;
     plaintext_out_size <= REG_COMB_plaintext_out_size;
     plaintext_remaining_out <= REG_COMB_plaintext_remaining_out;
     plaintext_out_expected <= REG_COMB_plaintext_out_expected;
     tag_match_checked <= REG_COMB_tag_match_checked;
 end if;
 end if;
end process;
-- Shared global regs
module_to_global.chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in when clk_en_internal='1' else chacha20poly1305_decrypt_axis_in;

end arch;
