-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 35
entity axis128_to_axis512_0CLK_c1f85885 is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 axis_in : in axis128_t_stream_t;
 axis_out_ready : in unsigned(0 downto 0);
 return_output : out axis128_to_axis512_t);
end axis128_to_axis512_0CLK_c1f85885;
architecture arch of axis128_to_axis512_0CLK_c1f85885 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal axis_in_reg : axis128_t_stream_t := axis128_t_stream_t_NULL;
signal axis_out_reg : axis512_t_stream_t := axis512_t_stream_t_NULL;
signal REG_COMB_axis_in_reg : axis128_t_stream_t;
signal REG_COMB_axis_out_reg : axis512_t_stream_t;

-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- BIN_OP_AND[axis_h_l377_c6_7d3c]
signal BIN_OP_AND_axis_h_l377_c6_7d3c_left : unsigned(0 downto 0);
signal BIN_OP_AND_axis_h_l377_c6_7d3c_right : unsigned(0 downto 0);
signal BIN_OP_AND_axis_h_l377_c6_7d3c_return_output : unsigned(0 downto 0);

-- axis_out_reg_data_tkeep_MUX[axis_h_l377_c3_425d]
signal axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_cond : unsigned(0 downto 0);
signal axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iftrue : uint1_t_64;
signal axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iffalse : uint1_t_64;
signal axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output : uint1_t_64;

-- axis_out_reg_data_tlast_MUX[axis_h_l377_c3_425d]
signal axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_cond : unsigned(0 downto 0);
signal axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iftrue : unsigned(0 downto 0);
signal axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iffalse : unsigned(0 downto 0);
signal axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output : unsigned(0 downto 0);

-- axis_out_reg_valid_MUX[axis_h_l377_c3_425d]
signal axis_out_reg_valid_MUX_axis_h_l377_c3_425d_cond : unsigned(0 downto 0);
signal axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iftrue : unsigned(0 downto 0);
signal axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iffalse : unsigned(0 downto 0);
signal axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output : unsigned(0 downto 0);

-- UNARY_OP_NOT[axis_h_l388_c28_5ae9]
signal UNARY_OP_NOT_axis_h_l388_c28_5ae9_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[axis_h_l389_c6_1ff2]
signal BIN_OP_AND_axis_h_l389_c6_1ff2_left : unsigned(0 downto 0);
signal BIN_OP_AND_axis_h_l389_c6_1ff2_right : unsigned(0 downto 0);
signal BIN_OP_AND_axis_h_l389_c6_1ff2_return_output : unsigned(0 downto 0);

-- axis_out_reg_MUX[axis_h_l389_c3_f755]
signal axis_out_reg_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
signal axis_out_reg_MUX_axis_h_l389_c3_f755_iftrue : axis512_t_stream_t;
signal axis_out_reg_MUX_axis_h_l389_c3_f755_iffalse : axis512_t_stream_t;
signal axis_out_reg_MUX_axis_h_l389_c3_f755_return_output : axis512_t_stream_t;

-- axis_in_reg_valid_MUX[axis_h_l389_c3_f755]
signal axis_in_reg_valid_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
signal axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iftrue : unsigned(0 downto 0);
signal axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iffalse : unsigned(0 downto 0);
signal axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output : unsigned(0 downto 0);

-- axis_in_reg_data_tkeep_MUX[axis_h_l389_c3_f755]
signal axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
signal axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iftrue : uint1_t_16;
signal axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iffalse : uint1_t_16;
signal axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output : uint1_t_16;

-- axis_in_reg_data_tlast_MUX[axis_h_l389_c3_f755]
signal axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
signal axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iftrue : unsigned(0 downto 0);
signal axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iffalse : unsigned(0 downto 0);
signal axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output : unsigned(0 downto 0);

-- axis512_to_axis128_array[axis_h_l393_c43_082a]
signal axis512_to_axis128_array_axis_h_l393_c43_082a_axis : axis512_t;
signal axis512_to_axis128_array_axis_h_l393_c43_082a_return_output : axis512_to_axis128_array_t;

-- axis_out_as_chunks_MUX[axis_h_l407_c5_498e]
signal axis_out_as_chunks_MUX_axis_h_l407_c5_498e_cond : unsigned(0 downto 0);
signal axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iftrue : axis128_t_stream_t_4;
signal axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iffalse : axis128_t_stream_t_4;
signal axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output : axis128_t_stream_t_4;

-- FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT[axis_h_l415_c13_96c5]
signal FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr : unsigned(0 downto 0);
signal FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX[axis_h_l415_c9_f506]
signal FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond : unsigned(0 downto 0);
signal FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue : axis128_t_stream_t_4;
signal FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse : axis128_t_stream_t_4;
signal FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;

-- FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT[axis_h_l415_c13_96c5]
signal FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr : unsigned(0 downto 0);
signal FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX[axis_h_l415_c9_f506]
signal FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond : unsigned(0 downto 0);
signal FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue : axis128_t_stream_t_4;
signal FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse : axis128_t_stream_t_4;
signal FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;

-- FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT[axis_h_l415_c13_96c5]
signal FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr : unsigned(0 downto 0);
signal FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output : unsigned(0 downto 0);

-- FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX[axis_h_l415_c9_f506]
signal FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond : unsigned(0 downto 0);
signal FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue : axis128_t_stream_t_4;
signal FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse : axis128_t_stream_t_4;
signal FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;

-- axis128_array_to_axis512[axis_h_l424_c25_67d5]
signal axis128_array_to_axis512_axis_h_l424_c25_67d5_axis_chunks : axis128_t_stream_t_4;
signal axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output : axis512_t;

-- UNARY_OP_NOT[axis_h_l432_c22_18b2]
signal UNARY_OP_NOT_axis_h_l432_c22_18b2_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[axis_h_l433_c6_0942]
signal BIN_OP_AND_axis_h_l433_c6_0942_left : unsigned(0 downto 0);
signal BIN_OP_AND_axis_h_l433_c6_0942_right : unsigned(0 downto 0);
signal BIN_OP_AND_axis_h_l433_c6_0942_return_output : unsigned(0 downto 0);

-- axis_in_reg_MUX[axis_h_l433_c3_0498]
signal axis_in_reg_MUX_axis_h_l433_c3_0498_cond : unsigned(0 downto 0);
signal axis_in_reg_MUX_axis_h_l433_c3_0498_iftrue : axis128_t_stream_t;
signal axis_in_reg_MUX_axis_h_l433_c3_0498_iffalse : axis128_t_stream_t;
signal axis_in_reg_MUX_axis_h_l433_c3_0498_return_output : axis128_t_stream_t;

function CONST_REF_RD_uint1_t_axis128_to_axis512_t_axis_out_valid_01c3( ref_toks_0 : axis512_t_stream_t) return unsigned is
 
  variable base : axis128_to_axis512_t; 
  variable return_output : unsigned(0 downto 0);
begin
      base.axis_out := ref_toks_0;

      return_output := base.axis_out.valid;
      return return_output; 
end function;

function CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_3b4a( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned) return uint1_t_64 is
 
  variable base : axis512_t_stream_t; 
  variable return_output : uint1_t_64;
begin
      base.data.tkeep(0) := ref_toks_0;
      base.data.tkeep(1) := ref_toks_1;
      base.data.tkeep(2) := ref_toks_2;
      base.data.tkeep(3) := ref_toks_3;
      base.data.tkeep(4) := ref_toks_4;
      base.data.tkeep(5) := ref_toks_5;
      base.data.tkeep(6) := ref_toks_6;
      base.data.tkeep(7) := ref_toks_7;
      base.data.tkeep(8) := ref_toks_8;
      base.data.tkeep(9) := ref_toks_9;
      base.data.tkeep(10) := ref_toks_10;
      base.data.tkeep(11) := ref_toks_11;
      base.data.tkeep(12) := ref_toks_12;
      base.data.tkeep(13) := ref_toks_13;
      base.data.tkeep(14) := ref_toks_14;
      base.data.tkeep(15) := ref_toks_15;
      base.data.tkeep(16) := ref_toks_16;
      base.data.tkeep(17) := ref_toks_17;
      base.data.tkeep(18) := ref_toks_18;
      base.data.tkeep(19) := ref_toks_19;
      base.data.tkeep(20) := ref_toks_20;
      base.data.tkeep(21) := ref_toks_21;
      base.data.tkeep(22) := ref_toks_22;
      base.data.tkeep(23) := ref_toks_23;
      base.data.tkeep(24) := ref_toks_24;
      base.data.tkeep(25) := ref_toks_25;
      base.data.tkeep(26) := ref_toks_26;
      base.data.tkeep(27) := ref_toks_27;
      base.data.tkeep(28) := ref_toks_28;
      base.data.tkeep(29) := ref_toks_29;
      base.data.tkeep(30) := ref_toks_30;
      base.data.tkeep(31) := ref_toks_31;
      base.data.tkeep(32) := ref_toks_32;
      base.data.tkeep(33) := ref_toks_33;
      base.data.tkeep(34) := ref_toks_34;
      base.data.tkeep(35) := ref_toks_35;
      base.data.tkeep(36) := ref_toks_36;
      base.data.tkeep(37) := ref_toks_37;
      base.data.tkeep(38) := ref_toks_38;
      base.data.tkeep(39) := ref_toks_39;
      base.data.tkeep(40) := ref_toks_40;
      base.data.tkeep(41) := ref_toks_41;
      base.data.tkeep(42) := ref_toks_42;
      base.data.tkeep(43) := ref_toks_43;
      base.data.tkeep(44) := ref_toks_44;
      base.data.tkeep(45) := ref_toks_45;
      base.data.tkeep(46) := ref_toks_46;
      base.data.tkeep(47) := ref_toks_47;
      base.data.tkeep(48) := ref_toks_48;
      base.data.tkeep(49) := ref_toks_49;
      base.data.tkeep(50) := ref_toks_50;
      base.data.tkeep(51) := ref_toks_51;
      base.data.tkeep(52) := ref_toks_52;
      base.data.tkeep(53) := ref_toks_53;
      base.data.tkeep(54) := ref_toks_54;
      base.data.tkeep(55) := ref_toks_55;
      base.data.tkeep(56) := ref_toks_56;
      base.data.tkeep(57) := ref_toks_57;
      base.data.tkeep(58) := ref_toks_58;
      base.data.tkeep(59) := ref_toks_59;
      base.data.tkeep(60) := ref_toks_60;
      base.data.tkeep(61) := ref_toks_61;
      base.data.tkeep(62) := ref_toks_62;
      base.data.tkeep(63) := ref_toks_63;

      return_output := base.data.tkeep;
      return return_output; 
end function;

function CONST_REF_RD_axis512_t_axis512_t_stream_t_data_699e( ref_toks_0 : axis512_t_stream_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : uint1_t_64) return axis512_t is
 
  variable base : axis512_t_stream_t; 
  variable return_output : axis512_t;
begin
      base := ref_toks_0;
      base.data.tlast := ref_toks_1;
      base.data.tkeep := ref_toks_2;

      return_output := base.data;
      return return_output; 
end function;

function CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_4e8d( ref_toks_0 : axis128_t_stream_t) return unsigned is
 
  variable base : axis128_t_stream_t_4; 
  variable return_output : unsigned(0 downto 0);
begin
      base(0) := ref_toks_0;

      return_output := base(0).valid;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346( ref_toks_0 : axis128_t_stream_t;
 ref_toks_1 : axis128_t_stream_t;
 ref_toks_2 : axis128_t_stream_t;
 ref_toks_3 : axis128_t_stream_t) return axis128_t_stream_t_4 is
 
  variable base : axis128_t_stream_t_4; 
  variable return_output : axis128_t_stream_t_4;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_42b0( ref_toks_0 : axis512_t;
 ref_toks_1 : unsigned) return axis512_t_stream_t is
 
  variable base : axis512_t_stream_t; 
  variable return_output : axis512_t_stream_t;
begin
      base.data := ref_toks_0;
      base.valid := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_6f11( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint1_t_16 is
 
  variable base : axis128_t_stream_t; 
  variable return_output : uint1_t_16;
begin
      base.data.tkeep(0) := ref_toks_0;
      base.data.tkeep(1) := ref_toks_1;
      base.data.tkeep(2) := ref_toks_2;
      base.data.tkeep(3) := ref_toks_3;
      base.data.tkeep(4) := ref_toks_4;
      base.data.tkeep(5) := ref_toks_5;
      base.data.tkeep(6) := ref_toks_6;
      base.data.tkeep(7) := ref_toks_7;
      base.data.tkeep(8) := ref_toks_8;
      base.data.tkeep(9) := ref_toks_9;
      base.data.tkeep(10) := ref_toks_10;
      base.data.tkeep(11) := ref_toks_11;
      base.data.tkeep(12) := ref_toks_12;
      base.data.tkeep(13) := ref_toks_13;
      base.data.tkeep(14) := ref_toks_14;
      base.data.tkeep(15) := ref_toks_15;

      return_output := base.data.tkeep;
      return return_output; 
end function;

function CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_4a8d( ref_toks_0 : axis512_t_stream_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : uint1_t_64) return axis512_t_stream_t is
 
  variable base : axis512_t_stream_t; 
  variable return_output : axis512_t_stream_t;
begin
      base := ref_toks_0;
      base.valid := ref_toks_1;
      base.data.tlast := ref_toks_2;
      base.data.tkeep := ref_toks_3;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_149c( ref_toks_0 : axis128_t_stream_t;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : uint1_t_16) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base := ref_toks_0;
      base.data.tlast := ref_toks_1;
      base.valid := ref_toks_2;
      base.data.tkeep := ref_toks_3;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_to_axis512_t_axis128_to_axis512_t_c1ed( ref_toks_0 : axis512_t_stream_t;
 ref_toks_1 : unsigned) return axis128_to_axis512_t is
 
  variable base : axis128_to_axis512_t; 
  variable return_output : axis128_to_axis512_t;
begin
      base.axis_out := ref_toks_0;
      base.axis_in_ready := ref_toks_1;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_AND_axis_h_l377_c6_7d3c : 0 clocks latency
BIN_OP_AND_axis_h_l377_c6_7d3c : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_axis_h_l377_c6_7d3c_left,
BIN_OP_AND_axis_h_l377_c6_7d3c_right,
BIN_OP_AND_axis_h_l377_c6_7d3c_return_output);

-- axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d : 0 clocks latency
axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d : entity work.MUX_uint1_t_uint1_t_64_uint1_t_64_0CLK_de264c78 port map (
axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_cond,
axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iftrue,
axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iffalse,
axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output);

-- axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d : 0 clocks latency
axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_cond,
axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iftrue,
axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iffalse,
axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output);

-- axis_out_reg_valid_MUX_axis_h_l377_c3_425d : 0 clocks latency
axis_out_reg_valid_MUX_axis_h_l377_c3_425d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
axis_out_reg_valid_MUX_axis_h_l377_c3_425d_cond,
axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iftrue,
axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iffalse,
axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output);

-- UNARY_OP_NOT_axis_h_l388_c28_5ae9 : 0 clocks latency
UNARY_OP_NOT_axis_h_l388_c28_5ae9 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_axis_h_l388_c28_5ae9_expr,
UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output);

-- BIN_OP_AND_axis_h_l389_c6_1ff2 : 0 clocks latency
BIN_OP_AND_axis_h_l389_c6_1ff2 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_axis_h_l389_c6_1ff2_left,
BIN_OP_AND_axis_h_l389_c6_1ff2_right,
BIN_OP_AND_axis_h_l389_c6_1ff2_return_output);

-- axis_out_reg_MUX_axis_h_l389_c3_f755 : 0 clocks latency
axis_out_reg_MUX_axis_h_l389_c3_f755 : entity work.MUX_uint1_t_axis512_t_stream_t_axis512_t_stream_t_0CLK_de264c78 port map (
axis_out_reg_MUX_axis_h_l389_c3_f755_cond,
axis_out_reg_MUX_axis_h_l389_c3_f755_iftrue,
axis_out_reg_MUX_axis_h_l389_c3_f755_iffalse,
axis_out_reg_MUX_axis_h_l389_c3_f755_return_output);

-- axis_in_reg_valid_MUX_axis_h_l389_c3_f755 : 0 clocks latency
axis_in_reg_valid_MUX_axis_h_l389_c3_f755 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
axis_in_reg_valid_MUX_axis_h_l389_c3_f755_cond,
axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iftrue,
axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iffalse,
axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output);

-- axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755 : 0 clocks latency
axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755 : entity work.MUX_uint1_t_uint1_t_16_uint1_t_16_0CLK_de264c78 port map (
axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_cond,
axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iftrue,
axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iffalse,
axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output);

-- axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755 : 0 clocks latency
axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_cond,
axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iftrue,
axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iffalse,
axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output);

-- axis512_to_axis128_array_axis_h_l393_c43_082a : 0 clocks latency
axis512_to_axis128_array_axis_h_l393_c43_082a : entity work.axis512_to_axis128_array_0CLK_4b8d8b28 port map (
axis512_to_axis128_array_axis_h_l393_c43_082a_axis,
axis512_to_axis128_array_axis_h_l393_c43_082a_return_output);

-- axis_out_as_chunks_MUX_axis_h_l407_c5_498e : 0 clocks latency
axis_out_as_chunks_MUX_axis_h_l407_c5_498e : entity work.MUX_uint1_t_axis128_t_stream_t_4_axis128_t_stream_t_4_0CLK_de264c78 port map (
axis_out_as_chunks_MUX_axis_h_l407_c5_498e_cond,
axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iftrue,
axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iffalse,
axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output);

-- FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5 : 0 clocks latency
FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr,
FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output);

-- FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506 : 0 clocks latency
FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506 : entity work.MUX_uint1_t_axis128_t_stream_t_4_axis128_t_stream_t_4_0CLK_de264c78 port map (
FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond,
FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue,
FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse,
FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output);

-- FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5 : 0 clocks latency
FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr,
FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output);

-- FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506 : 0 clocks latency
FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506 : entity work.MUX_uint1_t_axis128_t_stream_t_4_axis128_t_stream_t_4_0CLK_de264c78 port map (
FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond,
FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue,
FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse,
FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output);

-- FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5 : 0 clocks latency
FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr,
FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output);

-- FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506 : 0 clocks latency
FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506 : entity work.MUX_uint1_t_axis128_t_stream_t_4_axis128_t_stream_t_4_0CLK_de264c78 port map (
FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond,
FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue,
FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse,
FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output);

-- axis128_array_to_axis512_axis_h_l424_c25_67d5 : 0 clocks latency
axis128_array_to_axis512_axis_h_l424_c25_67d5 : entity work.axis128_array_to_axis512_0CLK_fcdf4ca0 port map (
axis128_array_to_axis512_axis_h_l424_c25_67d5_axis_chunks,
axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output);

-- UNARY_OP_NOT_axis_h_l432_c22_18b2 : 0 clocks latency
UNARY_OP_NOT_axis_h_l432_c22_18b2 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_axis_h_l432_c22_18b2_expr,
UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output);

-- BIN_OP_AND_axis_h_l433_c6_0942 : 0 clocks latency
BIN_OP_AND_axis_h_l433_c6_0942 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_axis_h_l433_c6_0942_left,
BIN_OP_AND_axis_h_l433_c6_0942_right,
BIN_OP_AND_axis_h_l433_c6_0942_return_output);

-- axis_in_reg_MUX_axis_h_l433_c3_0498 : 0 clocks latency
axis_in_reg_MUX_axis_h_l433_c3_0498 : entity work.MUX_uint1_t_axis128_t_stream_t_axis128_t_stream_t_0CLK_de264c78 port map (
axis_in_reg_MUX_axis_h_l433_c3_0498_cond,
axis_in_reg_MUX_axis_h_l433_c3_0498_iftrue,
axis_in_reg_MUX_axis_h_l433_c3_0498_iffalse,
axis_in_reg_MUX_axis_h_l433_c3_0498_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Inputs
 axis_in,
 axis_out_ready,
 -- Registers
 axis_in_reg,
 axis_out_reg,
 -- All submodule outputs
 BIN_OP_AND_axis_h_l377_c6_7d3c_return_output,
 axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output,
 axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output,
 axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output,
 UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output,
 BIN_OP_AND_axis_h_l389_c6_1ff2_return_output,
 axis_out_reg_MUX_axis_h_l389_c3_f755_return_output,
 axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output,
 axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output,
 axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output,
 axis512_to_axis128_array_axis_h_l393_c43_082a_return_output,
 axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output,
 FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output,
 FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output,
 FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output,
 FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output,
 FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output,
 FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output,
 axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output,
 UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output,
 BIN_OP_AND_axis_h_l433_c6_0942_return_output,
 axis_in_reg_MUX_axis_h_l433_c3_0498_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis128_to_axis512_t;
 variable VAR_axis_in : axis128_t_stream_t;
 variable VAR_axis_out_ready : unsigned(0 downto 0);
 variable VAR_IN_SIZE : unsigned(31 downto 0);
 variable VAR_OUT_SIZE : unsigned(31 downto 0);
 variable VAR_o : axis128_to_axis512_t;
 variable VAR_CONST_REF_RD_uint1_t_axis128_to_axis512_t_axis_out_valid_01c3_axis_h_l377_c6_dcc1_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_return_output : unsigned(0 downto 0);
 variable VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iftrue : uint1_t_64;
 variable VAR_axis_out_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_3b4a_axis_h_l377_c3_425d_return_output : uint1_t_64;
 variable VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iffalse : uint1_t_64;
 variable VAR_axis_out_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_d41d_axis_h_l377_c3_425d_return_output : uint1_t_64;
 variable VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output : uint1_t_64;
 variable VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_cond : unsigned(0 downto 0);
 variable VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iftrue : unsigned(0 downto 0);
 variable VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iffalse : unsigned(0 downto 0);
 variable VAR_axis_out_reg_data_tlast_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_data_tlast_d41d_axis_h_l377_c3_425d_return_output : unsigned(0 downto 0);
 variable VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output : unsigned(0 downto 0);
 variable VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_cond : unsigned(0 downto 0);
 variable VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iftrue : unsigned(0 downto 0);
 variable VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iffalse : unsigned(0 downto 0);
 variable VAR_axis_out_reg_valid_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_valid_d41d_axis_h_l377_c3_425d_return_output : unsigned(0 downto 0);
 variable VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output : unsigned(0 downto 0);
 variable VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_cond : unsigned(0 downto 0);
 variable VAR_ARRAY_SET_i : unsigned(31 downto 0);
 variable VAR_out_reg_ready : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_axis_h_l388_c28_5ae9_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_return_output : unsigned(0 downto 0);
 variable VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_iftrue : axis512_t_stream_t;
 variable VAR_axis_out_reg_TRUE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_42b0_axis_h_l389_c3_f755_return_output : axis512_t_stream_t;
 variable VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_iffalse : axis512_t_stream_t;
 variable VAR_axis_out_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_4a8d_axis_h_l389_c3_f755_return_output : axis512_t_stream_t;
 variable VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_return_output : axis512_t_stream_t;
 variable VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
 variable VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iftrue : unsigned(0 downto 0);
 variable VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iffalse : unsigned(0 downto 0);
 variable VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output : unsigned(0 downto 0);
 variable VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
 variable VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iftrue : uint1_t_16;
 variable VAR_axis_in_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_6f11_axis_h_l389_c3_f755_return_output : uint1_t_16;
 variable VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iffalse : uint1_t_16;
 variable VAR_axis_in_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_d41d_axis_h_l389_c3_f755_return_output : uint1_t_16;
 variable VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output : uint1_t_16;
 variable VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
 variable VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iftrue : unsigned(0 downto 0);
 variable VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iffalse : unsigned(0 downto 0);
 variable VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output : unsigned(0 downto 0);
 variable VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_cond : unsigned(0 downto 0);
 variable VAR_axis_out_as_chunks : axis128_t_stream_t_4;
 variable VAR_to_array : axis512_to_axis128_array_t;
 variable VAR_axis512_to_axis128_array_axis_h_l393_c43_082a_axis : axis512_t;
 variable VAR_CONST_REF_RD_axis512_t_axis512_t_stream_t_data_699e_axis_h_l393_c68_c2cd_return_output : axis512_t;
 variable VAR_axis512_to_axis128_array_axis_h_l393_c43_082a_return_output : axis512_to_axis128_array_t;
 variable VAR_CONST_REF_RD_axis128_t_stream_t_4_axis512_to_axis128_array_t_axis_chunks_d41d_axis_h_l394_c26_737a_return_output : axis128_t_stream_t_4;
 variable VAR_ARRAY_SHIFT_DOWN_i : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l398_c34_e128_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l398_c156_da7e_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l398_c34_e128_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l398_c156_da7e_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l398_c34_e128_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l398_c156_da7e_return_output : axis128_t_stream_t;
 variable VAR_last_cycle : unsigned(0 downto 0);
 variable VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iftrue : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;
 variable VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iffalse : axis128_t_stream_t_4;
 variable VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output : axis128_t_stream_t_4;
 variable VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_cond : unsigned(0 downto 0);
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_4e8d_axis_h_l415_c13_f2e6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond : unsigned(0 downto 0);
 variable VAR_NULL_CHUNK : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l415_c13_f2e6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l418_c162_f011_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l418_c162_f011_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l418_c162_f011_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l415_c13_f2e6_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse : axis128_t_stream_t_4;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l418_c162_f011_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l418_c162_f011_return_output : axis128_t_stream_t;
 variable VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l418_c162_f011_return_output : axis128_t_stream_t;
 variable VAR_axis128_array_to_axis512_axis_h_l424_c25_67d5_axis_chunks : axis128_t_stream_t_4;
 variable VAR_axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output : axis512_t;
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l427_c26_57f5_return_output : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l433_c6_d62c_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l433_c6_0942_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l433_c6_0942_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_axis_h_l433_c6_0942_return_output : unsigned(0 downto 0);
 variable VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_iftrue : axis128_t_stream_t;
 variable VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_iffalse : axis128_t_stream_t;
 variable VAR_axis_in_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_149c_axis_h_l433_c3_0498_return_output : axis128_t_stream_t;
 variable VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_return_output : axis128_t_stream_t;
 variable VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_axis128_to_axis512_t_axis128_to_axis512_t_c1ed_axis_h_l437_c10_3fe6_return_output : axis128_to_axis512_t;
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l389_DUPLICATE_773f_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_axis_h_l399_l389_DUPLICATE_dda9_return_output : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_l407_DUPLICATE_141b_return_output : axis128_t_stream_t_4;
 -- State registers comb logic variables
variable REG_VAR_axis_in_reg : axis128_t_stream_t;
variable REG_VAR_axis_out_reg : axis512_t_stream_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_axis_in_reg := axis_in_reg;
  REG_VAR_axis_out_reg := axis_out_reg;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iftrue := to_unsigned(0, 1);
     VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iftrue := to_unsigned(0, 1);
     VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iftrue := to_unsigned(0, 1);
     VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iftrue := to_unsigned(0, 1);
     -- axis_out_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_3b4a[axis_h_l377_c3_425d] LATENCY=0
     VAR_axis_out_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_3b4a_axis_h_l377_c3_425d_return_output := CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_3b4a(
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1));

     -- axis_in_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_6f11[axis_h_l389_c3_f755] LATENCY=0
     VAR_axis_in_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_6f11_axis_h_l389_c3_f755_return_output := CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_6f11(
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1),
     to_unsigned(0, 1));

     -- Submodule level 1
     VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iftrue := VAR_axis_in_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_6f11_axis_h_l389_c3_f755_return_output;
     VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iftrue := VAR_axis_out_reg_data_tkeep_TRUE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_3b4a_axis_h_l377_c3_425d_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;
     -- Mux in inputs
     VAR_axis_in := axis_in;
     VAR_axis_out_ready := axis_out_ready;

     -- Submodule level 0
     VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_iftrue := VAR_axis_in;
     VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_right := VAR_axis_out_ready;
     -- CONST_REF_RD_uint1_t_axis128_to_axis512_t_axis_out_valid_01c3[axis_h_l377_c6_dcc1] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_to_axis512_t_axis_out_valid_01c3_axis_h_l377_c6_dcc1_return_output := CONST_REF_RD_uint1_t_axis128_to_axis512_t_axis_out_valid_01c3(
     axis_out_reg);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l389_DUPLICATE_773f LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l389_DUPLICATE_773f_return_output := axis_in_reg.valid;

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_axis_h_l399_l389_DUPLICATE_dda9 LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_axis_h_l399_l389_DUPLICATE_dda9_return_output := axis_in_reg.data.tlast;

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d[axis_h_l433_c6_d62c] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l433_c6_d62c_return_output := VAR_axis_in.valid;

     -- axis_in_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_d41d[axis_h_l389_c3_f755] LATENCY=0
     VAR_axis_in_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_d41d_axis_h_l389_c3_f755_return_output := axis_in_reg.data.tkeep;

     -- axis_out_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_d41d[axis_h_l377_c3_425d] LATENCY=0
     VAR_axis_out_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_d41d_axis_h_l377_c3_425d_return_output := axis_out_reg.data.tkeep;

     -- axis_out_reg_valid_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_valid_d41d[axis_h_l377_c3_425d] LATENCY=0
     VAR_axis_out_reg_valid_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_valid_d41d_axis_h_l377_c3_425d_return_output := axis_out_reg.valid;

     -- axis_out_reg_data_tlast_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_data_tlast_d41d[axis_h_l377_c3_425d] LATENCY=0
     VAR_axis_out_reg_data_tlast_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_data_tlast_d41d_axis_h_l377_c3_425d_return_output := axis_out_reg.data.tlast;

     -- Submodule level 1
     VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iffalse := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_axis_h_l399_l389_DUPLICATE_dda9_return_output;
     VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_axis_h_l399_l389_DUPLICATE_dda9_return_output;
     VAR_BIN_OP_AND_axis_h_l433_c6_0942_left := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l433_c6_d62c_return_output;
     VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_left := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l389_DUPLICATE_773f_return_output;
     VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iffalse := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_axis_h_l389_DUPLICATE_773f_return_output;
     VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_left := VAR_CONST_REF_RD_uint1_t_axis128_to_axis512_t_axis_out_valid_01c3_axis_h_l377_c6_dcc1_return_output;
     VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iffalse := VAR_axis_in_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_16_axis128_t_stream_t_data_tkeep_d41d_axis_h_l389_c3_f755_return_output;
     VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iffalse := VAR_axis_out_reg_data_tkeep_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_64_axis512_t_stream_t_data_tkeep_d41d_axis_h_l377_c3_425d_return_output;
     VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iffalse := VAR_axis_out_reg_data_tlast_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_data_tlast_d41d_axis_h_l377_c3_425d_return_output;
     VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iffalse := VAR_axis_out_reg_valid_FALSE_INPUT_MUX_CONST_REF_RD_uint1_t_axis512_t_stream_t_valid_d41d_axis_h_l377_c3_425d_return_output;
     -- BIN_OP_AND[axis_h_l377_c6_7d3c] LATENCY=0
     -- Inputs
     BIN_OP_AND_axis_h_l377_c6_7d3c_left <= VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_left;
     BIN_OP_AND_axis_h_l377_c6_7d3c_right <= VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_right;
     -- Outputs
     VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_return_output := BIN_OP_AND_axis_h_l377_c6_7d3c_return_output;

     -- Submodule level 2
     VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_cond := VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_return_output;
     VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_cond := VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_return_output;
     VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_cond := VAR_BIN_OP_AND_axis_h_l377_c6_7d3c_return_output;
     -- axis_out_reg_data_tlast_MUX[axis_h_l377_c3_425d] LATENCY=0
     -- Inputs
     axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_cond <= VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_cond;
     axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iftrue <= VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iftrue;
     axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iffalse <= VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_iffalse;
     -- Outputs
     VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output := axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output;

     -- axis_out_reg_data_tkeep_MUX[axis_h_l377_c3_425d] LATENCY=0
     -- Inputs
     axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_cond <= VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_cond;
     axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iftrue <= VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iftrue;
     axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iffalse <= VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_iffalse;
     -- Outputs
     VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output := axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output;

     -- axis_out_reg_valid_MUX[axis_h_l377_c3_425d] LATENCY=0
     -- Inputs
     axis_out_reg_valid_MUX_axis_h_l377_c3_425d_cond <= VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_cond;
     axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iftrue <= VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iftrue;
     axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iffalse <= VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_iffalse;
     -- Outputs
     VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output := axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output;

     -- Submodule level 3
     VAR_UNARY_OP_NOT_axis_h_l388_c28_5ae9_expr := VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output;
     -- CONST_REF_RD_axis512_t_axis512_t_stream_t_data_699e[axis_h_l393_c68_c2cd] LATENCY=0
     VAR_CONST_REF_RD_axis512_t_axis512_t_stream_t_data_699e_axis_h_l393_c68_c2cd_return_output := CONST_REF_RD_axis512_t_axis512_t_stream_t_data_699e(
     axis_out_reg,
     VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output,
     VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output);

     -- UNARY_OP_NOT[axis_h_l388_c28_5ae9] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_axis_h_l388_c28_5ae9_expr <= VAR_UNARY_OP_NOT_axis_h_l388_c28_5ae9_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output := UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output;

     -- axis_out_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_4a8d[axis_h_l389_c3_f755] LATENCY=0
     VAR_axis_out_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_4a8d_axis_h_l389_c3_f755_return_output := CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_4a8d(
     axis_out_reg,
     VAR_axis_out_reg_valid_MUX_axis_h_l377_c3_425d_return_output,
     VAR_axis_out_reg_data_tlast_MUX_axis_h_l377_c3_425d_return_output,
     VAR_axis_out_reg_data_tkeep_MUX_axis_h_l377_c3_425d_return_output);

     -- Submodule level 4
     VAR_axis512_to_axis128_array_axis_h_l393_c43_082a_axis := VAR_CONST_REF_RD_axis512_t_axis512_t_stream_t_data_699e_axis_h_l393_c68_c2cd_return_output;
     VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_right := VAR_UNARY_OP_NOT_axis_h_l388_c28_5ae9_return_output;
     VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_iffalse := VAR_axis_out_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_4a8d_axis_h_l389_c3_f755_return_output;
     -- axis512_to_axis128_array[axis_h_l393_c43_082a] LATENCY=0
     -- Inputs
     axis512_to_axis128_array_axis_h_l393_c43_082a_axis <= VAR_axis512_to_axis128_array_axis_h_l393_c43_082a_axis;
     -- Outputs
     VAR_axis512_to_axis128_array_axis_h_l393_c43_082a_return_output := axis512_to_axis128_array_axis_h_l393_c43_082a_return_output;

     -- BIN_OP_AND[axis_h_l389_c6_1ff2] LATENCY=0
     -- Inputs
     BIN_OP_AND_axis_h_l389_c6_1ff2_left <= VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_left;
     BIN_OP_AND_axis_h_l389_c6_1ff2_right <= VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_right;
     -- Outputs
     VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_return_output := BIN_OP_AND_axis_h_l389_c6_1ff2_return_output;

     -- Submodule level 5
     VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_cond := VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_return_output;
     VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_cond := VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_return_output;
     VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_cond := VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_return_output;
     VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_cond := VAR_BIN_OP_AND_axis_h_l389_c6_1ff2_return_output;
     -- axis_in_reg_data_tlast_MUX[axis_h_l389_c3_f755] LATENCY=0
     -- Inputs
     axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_cond <= VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_cond;
     axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iftrue <= VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iftrue;
     axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iffalse <= VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_iffalse;
     -- Outputs
     VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output := axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output;

     -- CONST_REF_RD_axis128_t_stream_t_4_axis512_to_axis128_array_t_axis_chunks_d41d[axis_h_l394_c26_737a] LATENCY=0
     VAR_CONST_REF_RD_axis128_t_stream_t_4_axis512_to_axis128_array_t_axis_chunks_d41d_axis_h_l394_c26_737a_return_output := VAR_axis512_to_axis128_array_axis_h_l393_c43_082a_return_output.axis_chunks;

     -- axis_in_reg_valid_MUX[axis_h_l389_c3_f755] LATENCY=0
     -- Inputs
     axis_in_reg_valid_MUX_axis_h_l389_c3_f755_cond <= VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_cond;
     axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iftrue <= VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iftrue;
     axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iffalse <= VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_iffalse;
     -- Outputs
     VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output := axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output;

     -- axis_in_reg_data_tkeep_MUX[axis_h_l389_c3_f755] LATENCY=0
     -- Inputs
     axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_cond <= VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_cond;
     axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iftrue <= VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iftrue;
     axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iffalse <= VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_iffalse;
     -- Outputs
     VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output := axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output;

     -- Submodule level 6
     VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_expr := VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output;
     -- FOR_axis_h_l398_c34_e128_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d[axis_h_l398_c156_da7e] LATENCY=0
     VAR_FOR_axis_h_l398_c34_e128_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l398_c156_da7e_return_output := VAR_CONST_REF_RD_axis128_t_stream_t_4_axis512_to_axis128_array_t_axis_chunks_d41d_axis_h_l394_c26_737a_return_output(1);

     -- UNARY_OP_NOT[axis_h_l432_c22_18b2] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_axis_h_l432_c22_18b2_expr <= VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output := UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output;

     -- FOR_axis_h_l398_c34_e128_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d[axis_h_l398_c156_da7e] LATENCY=0
     VAR_FOR_axis_h_l398_c34_e128_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l398_c156_da7e_return_output := VAR_CONST_REF_RD_axis128_t_stream_t_4_axis512_to_axis128_array_t_axis_chunks_d41d_axis_h_l394_c26_737a_return_output(3);

     -- axis_in_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_149c[axis_h_l433_c3_0498] LATENCY=0
     VAR_axis_in_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_149c_axis_h_l433_c3_0498_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_149c(
     axis_in_reg,
     VAR_axis_in_reg_data_tlast_MUX_axis_h_l389_c3_f755_return_output,
     VAR_axis_in_reg_valid_MUX_axis_h_l389_c3_f755_return_output,
     VAR_axis_in_reg_data_tkeep_MUX_axis_h_l389_c3_f755_return_output);

     -- FOR_axis_h_l398_c34_e128_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d[axis_h_l398_c156_da7e] LATENCY=0
     VAR_FOR_axis_h_l398_c34_e128_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l398_c156_da7e_return_output := VAR_CONST_REF_RD_axis128_t_stream_t_4_axis512_to_axis128_array_t_axis_chunks_d41d_axis_h_l394_c26_737a_return_output(2);

     -- Submodule level 7
     VAR_BIN_OP_AND_axis_h_l433_c6_0942_right := VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output;
     VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_iffalse := VAR_axis_in_reg_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_149c_axis_h_l433_c3_0498_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346[axis_h_l415_c9_f506] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output := CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346(
     VAR_FOR_axis_h_l398_c34_e128_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l398_c156_da7e_return_output,
     VAR_FOR_axis_h_l398_c34_e128_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l398_c156_da7e_return_output,
     axis_in_reg,
     axis128_t_stream_t_NULL);

     -- CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_l407_DUPLICATE_141b LATENCY=0
     VAR_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_l407_DUPLICATE_141b_return_output := CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346(
     VAR_FOR_axis_h_l398_c34_e128_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l398_c156_da7e_return_output,
     VAR_FOR_axis_h_l398_c34_e128_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l398_c156_da7e_return_output,
     VAR_FOR_axis_h_l398_c34_e128_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l398_c156_da7e_return_output,
     axis_in_reg);

     -- BIN_OP_AND[axis_h_l433_c6_0942] LATENCY=0
     -- Inputs
     BIN_OP_AND_axis_h_l433_c6_0942_left <= VAR_BIN_OP_AND_axis_h_l433_c6_0942_left;
     BIN_OP_AND_axis_h_l433_c6_0942_right <= VAR_BIN_OP_AND_axis_h_l433_c6_0942_right;
     -- Outputs
     VAR_BIN_OP_AND_axis_h_l433_c6_0942_return_output := BIN_OP_AND_axis_h_l433_c6_0942_return_output;

     -- FOR_axis_h_l411_c7_ebdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_4e8d[axis_h_l415_c13_f2e6] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_4e8d_axis_h_l415_c13_f2e6_return_output := CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_4e8d(
     VAR_FOR_axis_h_l398_c34_e128_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l398_c156_da7e_return_output);

     -- CONST_REF_RD_axis128_to_axis512_t_axis128_to_axis512_t_c1ed[axis_h_l437_c10_3fe6] LATENCY=0
     VAR_CONST_REF_RD_axis128_to_axis512_t_axis128_to_axis512_t_c1ed_axis_h_l437_c10_3fe6_return_output := CONST_REF_RD_axis128_to_axis512_t_axis128_to_axis512_t_c1ed(
     axis_out_reg,
     VAR_UNARY_OP_NOT_axis_h_l432_c22_18b2_return_output);

     -- Submodule level 8
     VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_cond := VAR_BIN_OP_AND_axis_h_l433_c6_0942_return_output;
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse := VAR_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_l407_DUPLICATE_141b_return_output;
     VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iffalse := VAR_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_l407_DUPLICATE_141b_return_output;
     VAR_return_output := VAR_CONST_REF_RD_axis128_to_axis512_t_axis128_to_axis512_t_c1ed_axis_h_l437_c10_3fe6_return_output;
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_4e8d_axis_h_l415_c13_f2e6_return_output;
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT[axis_h_l415_c13_96c5] LATENCY=0
     -- Inputs
     FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr;
     -- Outputs
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output := FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output;

     -- axis_in_reg_MUX[axis_h_l433_c3_0498] LATENCY=0
     -- Inputs
     axis_in_reg_MUX_axis_h_l433_c3_0498_cond <= VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_cond;
     axis_in_reg_MUX_axis_h_l433_c3_0498_iftrue <= VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_iftrue;
     axis_in_reg_MUX_axis_h_l433_c3_0498_iffalse <= VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_iffalse;
     -- Outputs
     VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_return_output := axis_in_reg_MUX_axis_h_l433_c3_0498_return_output;

     -- Submodule level 9
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output;
     REG_VAR_axis_in_reg := VAR_axis_in_reg_MUX_axis_h_l433_c3_0498_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX[axis_h_l415_c9_f506] LATENCY=0
     -- Inputs
     FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond;
     FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue;
     FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse;
     -- Outputs
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output := FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output;

     -- Submodule level 10
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d[axis_h_l418_c162_f011] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l418_c162_f011_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(2);

     -- FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d[axis_h_l418_c162_f011] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l418_c162_f011_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(1);

     -- FOR_axis_h_l411_c7_ebdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d[axis_h_l415_c13_f2e6] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l415_c13_f2e6_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(0).valid;

     -- FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d[axis_h_l418_c162_f011] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l418_c162_f011_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_0_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(3);

     -- Submodule level 11
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l415_c13_f2e6_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346[axis_h_l415_c9_f506] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output := CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346(
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l418_c162_f011_return_output,
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l418_c162_f011_return_output,
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l418_c162_f011_return_output,
     axis128_t_stream_t_NULL);

     -- FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT[axis_h_l415_c13_96c5] LATENCY=0
     -- Inputs
     FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr;
     -- Outputs
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output := FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output;

     -- Submodule level 12
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output;
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX[axis_h_l415_c9_f506] LATENCY=0
     -- Inputs
     FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond;
     FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue;
     FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse;
     -- Outputs
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output := FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output;

     -- Submodule level 13
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d[axis_h_l415_c13_f2e6] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l415_c13_f2e6_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(0).valid;

     -- FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d[axis_h_l418_c162_f011] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l418_c162_f011_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(1);

     -- FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d[axis_h_l418_c162_f011] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l418_c162_f011_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(3);

     -- FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d[axis_h_l418_c162_f011] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l418_c162_f011_return_output := VAR_FOR_axis_h_l411_c7_ebdd_ITER_1_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output(2);

     -- Submodule level 14
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr := VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l415_c13_f2e6_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346[axis_h_l415_c9_f506] LATENCY=0
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output := CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346(
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_0_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_1_d41d_axis_h_l418_c162_f011_return_output,
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_1_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_2_d41d_axis_h_l418_c162_f011_return_output,
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_FOR_axis_h_l418_c40_10f7_ITER_2_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_4_3_d41d_axis_h_l418_c162_f011_return_output,
     axis128_t_stream_t_NULL);

     -- FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT[axis_h_l415_c13_96c5] LATENCY=0
     -- Inputs
     FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_expr;
     -- Outputs
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output := FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output;

     -- Submodule level 15
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond := VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_UNARY_OP_NOT_axis_h_l415_c13_96c5_return_output;
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue := VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_4_axis128_t_stream_t_4_2346_axis_h_l415_c9_f506_return_output;
     -- FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX[axis_h_l415_c9_f506] LATENCY=0
     -- Inputs
     FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_cond;
     FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iftrue;
     FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse <= VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_iffalse;
     -- Outputs
     VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output := FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output;

     -- Submodule level 16
     VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iftrue := VAR_FOR_axis_h_l411_c7_ebdd_ITER_2_axis_out_as_chunks_MUX_axis_h_l415_c9_f506_return_output;
     -- axis_out_as_chunks_MUX[axis_h_l407_c5_498e] LATENCY=0
     -- Inputs
     axis_out_as_chunks_MUX_axis_h_l407_c5_498e_cond <= VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_cond;
     axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iftrue <= VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iftrue;
     axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iffalse <= VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_iffalse;
     -- Outputs
     VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output := axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output;

     -- Submodule level 17
     VAR_axis128_array_to_axis512_axis_h_l424_c25_67d5_axis_chunks := VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output;
     -- axis128_array_to_axis512[axis_h_l424_c25_67d5] LATENCY=0
     -- Inputs
     axis128_array_to_axis512_axis_h_l424_c25_67d5_axis_chunks <= VAR_axis128_array_to_axis512_axis_h_l424_c25_67d5_axis_chunks;
     -- Outputs
     VAR_axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output := axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output;

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d[axis_h_l427_c26_57f5] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l427_c26_57f5_return_output := VAR_axis_out_as_chunks_MUX_axis_h_l407_c5_498e_return_output(0).valid;

     -- Submodule level 18
     -- axis_out_reg_TRUE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_42b0[axis_h_l389_c3_f755] LATENCY=0
     VAR_axis_out_reg_TRUE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_42b0_axis_h_l389_c3_f755_return_output := CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_42b0(
     VAR_axis128_array_to_axis512_axis_h_l424_c25_67d5_return_output,
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_4_0_valid_d41d_axis_h_l427_c26_57f5_return_output);

     -- Submodule level 19
     VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_iftrue := VAR_axis_out_reg_TRUE_INPUT_MUX_CONST_REF_RD_axis512_t_stream_t_axis512_t_stream_t_42b0_axis_h_l389_c3_f755_return_output;
     -- axis_out_reg_MUX[axis_h_l389_c3_f755] LATENCY=0
     -- Inputs
     axis_out_reg_MUX_axis_h_l389_c3_f755_cond <= VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_cond;
     axis_out_reg_MUX_axis_h_l389_c3_f755_iftrue <= VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_iftrue;
     axis_out_reg_MUX_axis_h_l389_c3_f755_iffalse <= VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_iffalse;
     -- Outputs
     VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_return_output := axis_out_reg_MUX_axis_h_l389_c3_f755_return_output;

     -- Submodule level 20
     REG_VAR_axis_out_reg := VAR_axis_out_reg_MUX_axis_h_l389_c3_f755_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_axis_in_reg <= REG_VAR_axis_in_reg;
REG_COMB_axis_out_reg <= REG_VAR_axis_out_reg;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     axis_in_reg <= REG_COMB_axis_in_reg;
     axis_out_reg <= REG_COMB_axis_out_reg;
 end if;
 end if;
end process;

end arch;
