mem['h0000] = 32'h00006517;
mem['h0001] = 32'h7E450513;
mem['h0002] = 32'h10000597;
mem['h0003] = 32'hFF858593;
mem['h0004] = 32'h10000617;
mem['h0005] = 32'hFF060613;
mem['h0006] = 32'h00C5DC63;
mem['h0007] = 32'h00052683;
mem['h0008] = 32'h00D5A023;
mem['h0009] = 32'h00450513;
mem['h000A] = 32'h00458593;
mem['h000B] = 32'hFEC5C8E3;
mem['h000C] = 32'h10000517;
mem['h000D] = 32'hFD050513;
mem['h000E] = 32'h10009597;
mem['h000F] = 32'hBF058593;
mem['h0010] = 32'h00B55863;
mem['h0011] = 32'h00052023;
mem['h0012] = 32'h00450513;
mem['h0013] = 32'hFEB54CE3;
mem['h0014] = 32'h10010117;
mem['h0015] = 32'hFB010113;
mem['h0016] = 32'h10000197;
mem['h0017] = 32'h7A818193;
mem['h0018] = 32'h00A54533;
mem['h0019] = 32'h00B5C5B3;
mem['h001A] = 32'h00C64633;
mem['h001B] = 32'h70D020EF;
mem['h001C] = 32'h0000006F;
mem['h001D] = 32'h00452783;
mem['h001E] = 32'h0087A783;
mem['h001F] = 32'h0007A783;
mem['h0020] = 32'h0007A783;
mem['h0021] = 32'hFE07C8E3;
mem['h0022] = 32'h00452783;
mem['h0023] = 32'h0087A783;
mem['h0024] = 32'h0007A783;
mem['h0025] = 32'h00B78023;
mem['h0026] = 32'h00008067;
mem['h0027] = 32'hFE010113;
mem['h0028] = 32'h00812C23;
mem['h0029] = 32'h01212823;
mem['h002A] = 32'hFFF60413;
mem['h002B] = 32'h00005937;
mem['h002C] = 32'h00912A23;
mem['h002D] = 32'h01312623;
mem['h002E] = 32'h00112E23;
mem['h002F] = 32'h00050493;
mem['h0030] = 32'h00058993;
mem['h0031] = 32'h00241413;
mem['h0032] = 32'h77090913;
mem['h0033] = 32'h0089D7B3;
mem['h0034] = 32'h00F7F793;
mem['h0035] = 32'h00F907B3;
mem['h0036] = 32'h0007C583;
mem['h0037] = 32'h00048513;
mem['h0038] = 32'hFFC40413;
mem['h0039] = 32'hF91FF0EF;
mem['h003A] = 32'hFE0452E3;
mem['h003B] = 32'h01C12083;
mem['h003C] = 32'h01812403;
mem['h003D] = 32'h01412483;
mem['h003E] = 32'h01012903;
mem['h003F] = 32'h00C12983;
mem['h0040] = 32'h02010113;
mem['h0041] = 32'h00008067;
mem['h0042] = 32'h0A058263;
mem['h0043] = 32'hFE010113;
mem['h0044] = 32'h00912A23;
mem['h0045] = 32'h00058493;
mem['h0046] = 32'h01212823;
mem['h0047] = 32'h00A00593;
mem['h0048] = 32'h00050913;
mem['h0049] = 32'h00048513;
mem['h004A] = 32'h00812C23;
mem['h004B] = 32'h00112E23;
mem['h004C] = 32'h01312623;
mem['h004D] = 32'h01412423;
mem['h004E] = 32'h00100413;
mem['h004F] = 32'h588050EF;
mem['h0050] = 32'h06857A63;
mem['h0051] = 32'h00900A13;
mem['h0052] = 32'h00040593;
mem['h0053] = 32'h00048513;
mem['h0054] = 32'h574050EF;
mem['h0055] = 32'h03050593;
mem['h0056] = 32'h0FF5F593;
mem['h0057] = 32'h00090513;
mem['h0058] = 32'hF15FF0EF;
mem['h0059] = 32'h00040593;
mem['h005A] = 32'h00048513;
mem['h005B] = 32'h5A0050EF;
mem['h005C] = 32'h00050493;
mem['h005D] = 32'h00A00593;
mem['h005E] = 32'h00040513;
mem['h005F] = 32'h00040993;
mem['h0060] = 32'h544050EF;
mem['h0061] = 32'h00050413;
mem['h0062] = 32'hFD3A60E3;
mem['h0063] = 32'h01C12083;
mem['h0064] = 32'h01812403;
mem['h0065] = 32'h01412483;
mem['h0066] = 32'h01012903;
mem['h0067] = 32'h00C12983;
mem['h0068] = 32'h00812A03;
mem['h0069] = 32'h02010113;
mem['h006A] = 32'h00008067;
mem['h006B] = 32'h03000593;
mem['h006C] = 32'hEC5FF06F;
mem['h006D] = 32'h00241793;
mem['h006E] = 32'h00878433;
mem['h006F] = 32'h00141413;
mem['h0070] = 32'hF81FF06F;
mem['h0071] = 32'hFF010113;
mem['h0072] = 32'h00812423;
mem['h0073] = 32'h00912223;
mem['h0074] = 32'h00112623;
mem['h0075] = 32'h00050493;
mem['h0076] = 32'h00058413;
mem['h0077] = 32'h00044583;
mem['h0078] = 32'h00059C63;
mem['h0079] = 32'h00C12083;
mem['h007A] = 32'h00812403;
mem['h007B] = 32'h00412483;
mem['h007C] = 32'h01010113;
mem['h007D] = 32'h00008067;
mem['h007E] = 32'h00048513;
mem['h007F] = 32'h00140413;
mem['h0080] = 32'hE75FF0EF;
mem['h0081] = 32'hFD9FF06F;
mem['h0082] = 32'hFF010113;
mem['h0083] = 32'h00112623;
mem['h0084] = 32'h00812423;
mem['h0085] = 32'h00912223;
mem['h0086] = 32'h00058493;
mem['h0087] = 32'h0005C583;
mem['h0088] = 32'h00050413;
mem['h0089] = 32'hEE5FF0EF;
mem['h008A] = 32'h00040513;
mem['h008B] = 32'h02E00593;
mem['h008C] = 32'hE45FF0EF;
mem['h008D] = 32'h0014C583;
mem['h008E] = 32'h00040513;
mem['h008F] = 32'hECDFF0EF;
mem['h0090] = 32'h00040513;
mem['h0091] = 32'h02E00593;
mem['h0092] = 32'hE2DFF0EF;
mem['h0093] = 32'h0024C583;
mem['h0094] = 32'h00040513;
mem['h0095] = 32'hEB5FF0EF;
mem['h0096] = 32'h00040513;
mem['h0097] = 32'h02E00593;
mem['h0098] = 32'hE15FF0EF;
mem['h0099] = 32'h00040513;
mem['h009A] = 32'h00812403;
mem['h009B] = 32'h0034C583;
mem['h009C] = 32'h00C12083;
mem['h009D] = 32'h00412483;
mem['h009E] = 32'h01010113;
mem['h009F] = 32'hE8DFF06F;
mem['h00A0] = 32'h00452783;
mem['h00A1] = 32'h0007A783;
mem['h00A2] = 32'h0007A783;
mem['h00A3] = 32'h0007A783;
mem['h00A4] = 32'h1407D863;
mem['h00A5] = 32'hFD010113;
mem['h00A6] = 32'h03212023;
mem['h00A7] = 32'h02112623;
mem['h00A8] = 32'h02812423;
mem['h00A9] = 32'h02912223;
mem['h00AA] = 32'h01312E23;
mem['h00AB] = 32'h01412C23;
mem['h00AC] = 32'h01512A23;
mem['h00AD] = 32'h01612823;
mem['h00AE] = 32'h01712623;
mem['h00AF] = 32'h0FF7F713;
mem['h00B0] = 32'h01200693;
mem['h00B1] = 32'h00050913;
mem['h00B2] = 32'h00000513;
mem['h00B3] = 32'h0AD70263;
mem['h00B4] = 32'h00058493;
mem['h00B5] = 32'h0FF7F593;
mem['h00B6] = 32'h00B48023;
mem['h00B7] = 32'h00A00793;
mem['h00B8] = 32'h0AF58E63;
mem['h00B9] = 32'h00D00793;
mem['h00BA] = 32'h00000413;
mem['h00BB] = 32'h0AF58E63;
mem['h00BC] = 32'h00800A13;
mem['h00BD] = 32'h07F00A93;
mem['h00BE] = 32'h01F00993;
mem['h00BF] = 32'h00A00B13;
mem['h00C0] = 32'h00D00B93;
mem['h00C1] = 32'h01458463;
mem['h00C2] = 32'h0D559263;
mem['h00C3] = 32'h02805863;
mem['h00C4] = 32'h00800593;
mem['h00C5] = 32'h00090513;
mem['h00C6] = 32'hD5DFF0EF;
mem['h00C7] = 32'h02000593;
mem['h00C8] = 32'h00090513;
mem['h00C9] = 32'hD51FF0EF;
mem['h00CA] = 32'h00800593;
mem['h00CB] = 32'h00090513;
mem['h00CC] = 32'hFFF48493;
mem['h00CD] = 32'hFFF40413;
mem['h00CE] = 32'hD3DFF0EF;
mem['h00CF] = 32'h00492783;
mem['h00D0] = 32'h0007A783;
mem['h00D1] = 32'h0007A783;
mem['h00D2] = 32'h0007A783;
mem['h00D3] = 32'hFE07D8E3;
mem['h00D4] = 32'h01340C63;
mem['h00D5] = 32'h0FF7F593;
mem['h00D6] = 32'h00B48023;
mem['h00D7] = 32'h05659463;
mem['h00D8] = 32'h00148493;
mem['h00D9] = 32'h00140413;
mem['h00DA] = 32'h00048023;
mem['h00DB] = 32'h0FF47513;
mem['h00DC] = 32'h02C12083;
mem['h00DD] = 32'h02812403;
mem['h00DE] = 32'h02412483;
mem['h00DF] = 32'h02012903;
mem['h00E0] = 32'h01C12983;
mem['h00E1] = 32'h01812A03;
mem['h00E2] = 32'h01412A83;
mem['h00E3] = 32'h01012B03;
mem['h00E4] = 32'h00C12B83;
mem['h00E5] = 32'h03010113;
mem['h00E6] = 32'h00008067;
mem['h00E7] = 32'h00000413;
mem['h00E8] = 32'hFC1FF06F;
mem['h00E9] = 32'hF77590E3;
mem['h00EA] = 32'h00D00593;
mem['h00EB] = 32'h00090513;
mem['h00EC] = 32'hCC5FF0EF;
mem['h00ED] = 32'h00A00593;
mem['h00EE] = 32'h00090513;
mem['h00EF] = 32'hCB9FF0EF;
mem['h00F0] = 32'h00A00793;
mem['h00F1] = 32'h00F48023;
mem['h00F2] = 32'hF99FF06F;
mem['h00F3] = 32'h00090513;
mem['h00F4] = 32'hCA5FF0EF;
mem['h00F5] = 32'h00148493;
mem['h00F6] = 32'h00140413;
mem['h00F7] = 32'hF61FF06F;
mem['h00F8] = 32'h00000513;
mem['h00F9] = 32'h00008067;
mem['h00FA] = 32'h00100613;
mem['h00FB] = 32'h00010837;
mem['h00FC] = 32'h00050693;
mem['h00FD] = 32'h00000793;
mem['h00FE] = 32'h40A60633;
mem['h00FF] = 32'hFFF80893;
mem['h0100] = 32'h00D60733;
mem['h0101] = 32'h04B76063;
mem['h0102] = 32'hFFE5F713;
mem['h0103] = 32'h02B77463;
mem['h0104] = 32'h00E50533;
mem['h0105] = 32'h00054703;
mem['h0106] = 32'h00871713;
mem['h0107] = 32'h00E787B3;
mem['h0108] = 32'h00010737;
mem['h0109] = 32'h00E7E863;
mem['h010A] = 32'h01079793;
mem['h010B] = 32'h0107D793;
mem['h010C] = 32'h00178793;
mem['h010D] = 32'hFFF7C513;
mem['h010E] = 32'h01051513;
mem['h010F] = 32'h01055513;
mem['h0110] = 32'h00008067;
mem['h0111] = 32'h0006C703;
mem['h0112] = 32'h0016C303;
mem['h0113] = 32'h00871713;
mem['h0114] = 32'h00676733;
mem['h0115] = 32'h01071713;
mem['h0116] = 32'h01075713;
mem['h0117] = 32'h00E787B3;
mem['h0118] = 32'h0107E663;
mem['h0119] = 32'h0117F7B3;
mem['h011A] = 32'h00178793;
mem['h011B] = 32'h00268693;
mem['h011C] = 32'hF91FF06F;
mem['h011D] = 32'h00000713;
mem['h011E] = 32'h00C71663;
mem['h011F] = 32'h00000513;
mem['h0120] = 32'h00008067;
mem['h0121] = 32'h00E507B3;
mem['h0122] = 32'h00E586B3;
mem['h0123] = 32'h0007C783;
mem['h0124] = 32'h0006C683;
mem['h0125] = 32'h00D78663;
mem['h0126] = 32'h40D78533;
mem['h0127] = 32'h00008067;
mem['h0128] = 32'h00170713;
mem['h0129] = 32'hFD5FF06F;
mem['h012A] = 32'h00050793;
mem['h012B] = 32'h00000513;
mem['h012C] = 32'h00A78733;
mem['h012D] = 32'h00074703;
mem['h012E] = 32'h00071463;
mem['h012F] = 32'h00008067;
mem['h0130] = 32'h00150513;
mem['h0131] = 32'hFEDFF06F;
mem['h0132] = 32'hFE010113;
mem['h0133] = 32'h00812C23;
mem['h0134] = 32'h00112E23;
mem['h0135] = 32'h00050413;
mem['h0136] = 32'h00B12623;
mem['h0137] = 32'hFCDFF0EF;
mem['h0138] = 32'h00050613;
mem['h0139] = 32'h00040513;
mem['h013A] = 32'h01812403;
mem['h013B] = 32'h00C12583;
mem['h013C] = 32'h01C12083;
mem['h013D] = 32'h02010113;
mem['h013E] = 32'hF7DFF06F;
mem['h013F] = 32'h00050813;
mem['h0140] = 32'h00054503;
mem['h0141] = 32'h00A00793;
mem['h0142] = 32'h06F50463;
mem['h0143] = 32'h06050463;
mem['h0144] = 32'h00000713;
mem['h0145] = 32'h00A00893;
mem['h0146] = 32'h00900313;
mem['h0147] = 32'h00084503;
mem['h0148] = 32'h01151863;
mem['h0149] = 32'h00000513;
mem['h014A] = 32'h02C77A63;
mem['h014B] = 32'h00008067;
mem['h014C] = 32'hFE050AE3;
mem['h014D] = 32'hFD050793;
mem['h014E] = 32'h0FF7F793;
mem['h014F] = 32'h02F36A63;
mem['h0150] = 32'h00271793;
mem['h0151] = 32'h00E787B3;
mem['h0152] = 32'h00179793;
mem['h0153] = 32'hFD078793;
mem['h0154] = 32'h00F50733;
mem['h0155] = 32'h00180813;
mem['h0156] = 32'hFC5FF06F;
mem['h0157] = 32'h00000513;
mem['h0158] = 32'h00E6EA63;
mem['h0159] = 32'h00E5A023;
mem['h015A] = 32'h00100513;
mem['h015B] = 32'h00008067;
mem['h015C] = 32'h00000513;
mem['h015D] = 32'h00008067;
mem['h015E] = 32'h0005A703;
mem['h015F] = 32'h00052783;
mem['h0160] = 32'h00E787B3;
mem['h0161] = 32'h00F52023;
mem['h0162] = 32'h0006A703;
mem['h0163] = 32'h00E7C7B3;
mem['h0164] = 32'h01079713;
mem['h0165] = 32'h0107D793;
mem['h0166] = 32'h00E7E7B3;
mem['h0167] = 32'h00F6A023;
mem['h0168] = 32'h00062703;
mem['h0169] = 32'h00E787B3;
mem['h016A] = 32'h00F62023;
mem['h016B] = 32'h0005A703;
mem['h016C] = 32'h00E7C7B3;
mem['h016D] = 32'h00C79713;
mem['h016E] = 32'h0147D793;
mem['h016F] = 32'h00E7E7B3;
mem['h0170] = 32'h00F5A023;
mem['h0171] = 32'h00052703;
mem['h0172] = 32'h00E787B3;
mem['h0173] = 32'h00F52023;
mem['h0174] = 32'h0006A703;
mem['h0175] = 32'h00E7C7B3;
mem['h0176] = 32'h00879713;
mem['h0177] = 32'h0187D793;
mem['h0178] = 32'h00E7E7B3;
mem['h0179] = 32'h00F6A023;
mem['h017A] = 32'h00062703;
mem['h017B] = 32'h00E787B3;
mem['h017C] = 32'h00F62023;
mem['h017D] = 32'h0005A703;
mem['h017E] = 32'h00E7C7B3;
mem['h017F] = 32'h00779713;
mem['h0180] = 32'h0197D793;
mem['h0181] = 32'h00F767B3;
mem['h0182] = 32'h00F5A023;
mem['h0183] = 32'h00008067;
mem['h0184] = 32'h00000693;
mem['h0185] = 32'h00000713;
mem['h0186] = 32'h02800E93;
mem['h0187] = 32'h00D587B3;
mem['h0188] = 32'h00D60833;
mem['h0189] = 32'h0007A303;
mem['h018A] = 32'h0047A883;
mem['h018B] = 32'h00082783;
mem['h018C] = 32'h00482803;
mem['h018D] = 32'h00F307B3;
mem['h018E] = 32'h0067BE33;
mem['h018F] = 32'h01088833;
mem['h0190] = 32'h010E0E33;
mem['h0191] = 32'h00E78833;
mem['h0192] = 32'h00F837B3;
mem['h0193] = 32'h01C787B3;
mem['h0194] = 32'h0317E063;
mem['h0195] = 32'h00F89463;
mem['h0196] = 32'h00686C63;
mem['h0197] = 32'h01031663;
mem['h0198] = 32'h00177713;
mem['h0199] = 32'h00F88863;
mem['h019A] = 32'h00000713;
mem['h019B] = 32'h0080006F;
mem['h019C] = 32'h00100713;
mem['h019D] = 32'h00D508B3;
mem['h019E] = 32'h0108A023;
mem['h019F] = 32'h00F8A223;
mem['h01A0] = 32'h00868693;
mem['h01A1] = 32'hF9D69CE3;
mem['h01A2] = 32'h00008067;
mem['h01A3] = 32'h0085D793;
mem['h01A4] = 32'h00B50023;
mem['h01A5] = 32'h00F500A3;
mem['h01A6] = 32'h0105D793;
mem['h01A7] = 32'h0185D593;
mem['h01A8] = 32'h00F50123;
mem['h01A9] = 32'h00B501A3;
mem['h01AA] = 32'h00050223;
mem['h01AB] = 32'h000502A3;
mem['h01AC] = 32'h00050323;
mem['h01AD] = 32'h000503A3;
mem['h01AE] = 32'h00008067;
mem['h01AF] = 32'hFD010113;
mem['h01B0] = 32'h02812423;
mem['h01B1] = 32'h01612823;
mem['h01B2] = 32'h01712623;
mem['h01B3] = 32'h01812423;
mem['h01B4] = 32'h01912223;
mem['h01B5] = 32'h01A12023;
mem['h01B6] = 32'h02112623;
mem['h01B7] = 32'h02912223;
mem['h01B8] = 32'h03212023;
mem['h01B9] = 32'h01312E23;
mem['h01BA] = 32'h01412C23;
mem['h01BB] = 32'h01512A23;
mem['h01BC] = 32'h00050B93;
mem['h01BD] = 32'h00050413;
mem['h01BE] = 32'h00000B13;
mem['h01BF] = 32'h00010D37;
mem['h01C0] = 32'hFFFF0CB7;
mem['h01C1] = 32'h01000C13;
mem['h01C2] = 32'h00042903;
mem['h01C3] = 32'h00442783;
mem['h01C4] = 32'h000B0713;
mem['h01C5] = 32'h01A904B3;
mem['h01C6] = 32'h0124B933;
mem['h01C7] = 32'h00F90933;
mem['h01C8] = 32'h00942023;
mem['h01C9] = 32'h01242223;
mem['h01CA] = 32'h00F72793;
mem['h01CB] = 32'h001B0B13;
mem['h01CC] = 32'h00000993;
mem['h01CD] = 32'h00078463;
mem['h01CE] = 32'h000B0993;
mem['h01CF] = 32'h01091693;
mem['h01D0] = 32'h0104D793;
mem['h01D1] = 32'h00F6E7B3;
mem['h01D2] = 32'h00399993;
mem['h01D3] = 32'h41095A93;
mem['h01D4] = 32'hFFF78A13;
mem['h01D5] = 32'hFF170713;
mem['h01D6] = 32'h0017B793;
mem['h01D7] = 32'h013B89B3;
mem['h01D8] = 32'h40FA8AB3;
mem['h01D9] = 32'h0A071663;
mem['h01DA] = 32'h000A0513;
mem['h01DB] = 32'h000A8593;
mem['h01DC] = 32'h00000693;
mem['h01DD] = 32'h02500613;
mem['h01DE] = 32'h6B9040EF;
mem['h01DF] = 32'h0009A703;
mem['h01E0] = 32'h0049A683;
mem['h01E1] = 32'h01450A33;
mem['h01E2] = 32'h00AA37B3;
mem['h01E3] = 32'h015585B3;
mem['h01E4] = 32'h01470A33;
mem['h01E5] = 32'h00B787B3;
mem['h01E6] = 32'h00F687B3;
mem['h01E7] = 32'h00EA3733;
mem['h01E8] = 32'h00F70733;
mem['h01E9] = 32'h0149A023;
mem['h01EA] = 32'h00E9A223;
mem['h01EB] = 32'h00042703;
mem['h01EC] = 32'h00442783;
mem['h01ED] = 32'h009CF4B3;
mem['h01EE] = 32'h409704B3;
mem['h01EF] = 32'h00973733;
mem['h01F0] = 32'h412787B3;
mem['h01F1] = 32'h40E787B3;
mem['h01F2] = 32'h00942023;
mem['h01F3] = 32'h00F42223;
mem['h01F4] = 32'h00840413;
mem['h01F5] = 32'hF38B1AE3;
mem['h01F6] = 32'h02C12083;
mem['h01F7] = 32'h02812403;
mem['h01F8] = 32'h02412483;
mem['h01F9] = 32'h02012903;
mem['h01FA] = 32'h01C12983;
mem['h01FB] = 32'h01812A03;
mem['h01FC] = 32'h01412A83;
mem['h01FD] = 32'h01012B03;
mem['h01FE] = 32'h00C12B83;
mem['h01FF] = 32'h00812C03;
mem['h0200] = 32'h00412C83;
mem['h0201] = 32'h00012D03;
mem['h0202] = 32'h03010113;
mem['h0203] = 32'h00008067;
mem['h0204] = 32'h00000513;
mem['h0205] = 32'h00000593;
mem['h0206] = 32'hF59FF06F;
mem['h0207] = 32'hFE010113;
mem['h0208] = 32'h00812C23;
mem['h0209] = 32'h00912A23;
mem['h020A] = 32'h01212823;
mem['h020B] = 32'h01312623;
mem['h020C] = 32'h01412423;
mem['h020D] = 32'h01512223;
mem['h020E] = 32'h00112E23;
mem['h020F] = 32'h00060913;
mem['h0210] = 32'h00050493;
mem['h0211] = 32'h00058413;
mem['h0212] = 32'h08058A13;
mem['h0213] = 32'h00167A93;
mem['h0214] = 32'h41F65993;
mem['h0215] = 32'h0004A503;
mem['h0216] = 32'h0044A583;
mem['h0217] = 32'h00042703;
mem['h0218] = 32'h00442783;
mem['h0219] = 32'h060A8863;
mem['h021A] = 32'h00070693;
mem['h021B] = 32'h00078613;
mem['h021C] = 32'h00D4A023;
mem['h021D] = 32'h00C4A223;
mem['h021E] = 32'h00F5C5B3;
mem['h021F] = 32'h00090613;
mem['h0220] = 32'h00098693;
mem['h0221] = 32'h00E54533;
mem['h0222] = 32'h5A9040EF;
mem['h0223] = 32'h00042783;
mem['h0224] = 32'h00840413;
mem['h0225] = 32'h00848493;
mem['h0226] = 32'h00A7C533;
mem['h0227] = 32'hFFC42783;
mem['h0228] = 32'hFEA42C23;
mem['h0229] = 32'h00B7C7B3;
mem['h022A] = 32'hFEF42E23;
mem['h022B] = 32'hFB4414E3;
mem['h022C] = 32'h01C12083;
mem['h022D] = 32'h01812403;
mem['h022E] = 32'h01412483;
mem['h022F] = 32'h01012903;
mem['h0230] = 32'h00C12983;
mem['h0231] = 32'h00812A03;
mem['h0232] = 32'h00412A83;
mem['h0233] = 32'h02010113;
mem['h0234] = 32'h00008067;
mem['h0235] = 32'h00050693;
mem['h0236] = 32'h00058613;
mem['h0237] = 32'hF95FF06F;
mem['h0238] = 32'h00000793;
mem['h0239] = 32'h08000E13;
mem['h023A] = 32'h00F586B3;
mem['h023B] = 32'h00F60333;
mem['h023C] = 32'h0006A703;
mem['h023D] = 32'h0046A803;
mem['h023E] = 32'h00032683;
mem['h023F] = 32'h00432303;
mem['h0240] = 32'h00F508B3;
mem['h0241] = 32'h00D706B3;
mem['h0242] = 32'h00E6B733;
mem['h0243] = 32'h00680833;
mem['h0244] = 32'h01070733;
mem['h0245] = 32'h00D8A023;
mem['h0246] = 32'h00E8A223;
mem['h0247] = 32'h00878793;
mem['h0248] = 32'hFDC794E3;
mem['h0249] = 32'h00008067;
mem['h024A] = 32'h00000793;
mem['h024B] = 32'h08000E13;
mem['h024C] = 32'h00F58733;
mem['h024D] = 32'h00F60333;
mem['h024E] = 32'h00072803;
mem['h024F] = 32'h00032683;
mem['h0250] = 32'h00472703;
mem['h0251] = 32'h00432303;
mem['h0252] = 32'h40D806B3;
mem['h0253] = 32'h00D83833;
mem['h0254] = 32'h40670733;
mem['h0255] = 32'h00F508B3;
mem['h0256] = 32'h41070733;
mem['h0257] = 32'h00D8A023;
mem['h0258] = 32'h00E8A223;
mem['h0259] = 32'h00878793;
mem['h025A] = 32'hFDC794E3;
mem['h025B] = 32'h00008067;
mem['h025C] = 32'hEC010113;
mem['h025D] = 32'h12812C23;
mem['h025E] = 32'h01810413;
mem['h025F] = 32'h13412623;
mem['h0260] = 32'h13512423;
mem['h0261] = 32'h13712023;
mem['h0262] = 32'h11A12A23;
mem['h0263] = 32'h12112E23;
mem['h0264] = 32'h12912A23;
mem['h0265] = 32'h13212823;
mem['h0266] = 32'h13612223;
mem['h0267] = 32'h11812E23;
mem['h0268] = 32'h11912C23;
mem['h0269] = 32'h11B12823;
mem['h026A] = 32'h00050A13;
mem['h026B] = 32'h00058D13;
mem['h026C] = 32'h00060B93;
mem['h026D] = 32'h00040793;
mem['h026E] = 32'h00040A93;
mem['h026F] = 32'h00000713;
mem['h0270] = 32'h00000693;
mem['h0271] = 32'h00E7A223;
mem['h0272] = 32'h00D7A023;
mem['h0273] = 32'h11010713;
mem['h0274] = 32'h00878793;
mem['h0275] = 32'hFEE794E3;
mem['h0276] = 32'h00040C93;
mem['h0277] = 32'h00000C13;
mem['h0278] = 32'h080B8D93;
mem['h0279] = 32'h01000913;
mem['h027A] = 32'h003C1793;
mem['h027B] = 32'h00FD07B3;
mem['h027C] = 32'h0047A803;
mem['h027D] = 32'h0007A783;
mem['h027E] = 32'h000B8B13;
mem['h027F] = 32'h01012623;
mem['h0280] = 32'h00F12423;
mem['h0281] = 32'h000C8493;
mem['h0282] = 32'h000B2603;
mem['h0283] = 32'h004B2683;
mem['h0284] = 32'h00812503;
mem['h0285] = 32'h00C12583;
mem['h0286] = 32'h008B0B13;
mem['h0287] = 32'h00848493;
mem['h0288] = 32'h411040EF;
mem['h0289] = 32'hFF84A783;
mem['h028A] = 32'hFFC4A703;
mem['h028B] = 32'h00A78533;
mem['h028C] = 32'h00F537B3;
mem['h028D] = 32'h00B70733;
mem['h028E] = 32'h00E787B3;
mem['h028F] = 32'hFEA4AC23;
mem['h0290] = 32'hFEF4AE23;
mem['h0291] = 32'hFDBB12E3;
mem['h0292] = 32'h001C0C13;
mem['h0293] = 32'h008C8C93;
mem['h0294] = 32'hF92C1CE3;
mem['h0295] = 32'h07840493;
mem['h0296] = 32'h08042503;
mem['h0297] = 32'h08442583;
mem['h0298] = 32'h02600613;
mem['h0299] = 32'h00000693;
mem['h029A] = 32'h3C9040EF;
mem['h029B] = 32'h00042783;
mem['h029C] = 32'h00442703;
mem['h029D] = 32'h00840413;
mem['h029E] = 32'h00A78533;
mem['h029F] = 32'h00F537B3;
mem['h02A0] = 32'h00B70733;
mem['h02A1] = 32'h00E787B3;
mem['h02A2] = 32'hFEA42C23;
mem['h02A3] = 32'hFEF42E23;
mem['h02A4] = 32'hFC8494E3;
mem['h02A5] = 32'h00000793;
mem['h02A6] = 32'h08000713;
mem['h02A7] = 32'h00FA8633;
mem['h02A8] = 32'h00062503;
mem['h02A9] = 32'h00462583;
mem['h02AA] = 32'h00FA06B3;
mem['h02AB] = 32'h00A6A023;
mem['h02AC] = 32'h00B6A223;
mem['h02AD] = 32'h00878793;
mem['h02AE] = 32'hFEE792E3;
mem['h02AF] = 32'h000A0513;
mem['h02B0] = 32'hBFDFF0EF;
mem['h02B1] = 32'h13812403;
mem['h02B2] = 32'h13C12083;
mem['h02B3] = 32'h13412483;
mem['h02B4] = 32'h13012903;
mem['h02B5] = 32'h12812A83;
mem['h02B6] = 32'h12412B03;
mem['h02B7] = 32'h12012B83;
mem['h02B8] = 32'h11C12C03;
mem['h02B9] = 32'h11812C83;
mem['h02BA] = 32'h11412D03;
mem['h02BB] = 32'h11012D83;
mem['h02BC] = 32'h000A0513;
mem['h02BD] = 32'h12C12A03;
mem['h02BE] = 32'h14010113;
mem['h02BF] = 32'hBC1FF06F;
mem['h02C0] = 32'hEC010113;
mem['h02C1] = 32'h13212823;
mem['h02C2] = 32'h00058913;
mem['h02C3] = 32'h000065B7;
mem['h02C4] = 32'h12812C23;
mem['h02C5] = 32'h12912A23;
mem['h02C6] = 32'h00050413;
mem['h02C7] = 32'h63058493;
mem['h02C8] = 32'h0A000613;
mem['h02C9] = 32'h63058593;
mem['h02CA] = 32'h08010513;
mem['h02CB] = 32'h12112E23;
mem['h02CC] = 32'h13312623;
mem['h02CD] = 32'h13412423;
mem['h02CE] = 32'h13512223;
mem['h02CF] = 32'h13612023;
mem['h02D0] = 32'h2C1010EF;
mem['h02D1] = 32'h04040E13;
mem['h02D2] = 32'h04010E93;
mem['h02D3] = 32'h0A048793;
mem['h02D4] = 32'h00040693;
mem['h02D5] = 32'h06040F13;
mem['h02D6] = 32'h000E8613;
mem['h02D7] = 32'h000E0713;
mem['h02D8] = 32'h00072583;
mem['h02D9] = 32'h00470713;
mem['h02DA] = 32'h00460613;
mem['h02DB] = 32'hFEB62E23;
mem['h02DC] = 32'h0007A583;
mem['h02DD] = 32'h00478793;
mem['h02DE] = 32'h00B62E23;
mem['h02DF] = 32'hFEEF12E3;
mem['h02E0] = 32'h06042783;
mem['h02E1] = 32'h07012883;
mem['h02E2] = 32'h06442703;
mem['h02E3] = 32'h00F8C8B3;
mem['h02E4] = 32'h07412783;
mem['h02E5] = 32'h00E7C7B3;
mem['h02E6] = 32'h00090863;
mem['h02E7] = 32'h07812703;
mem['h02E8] = 32'hFFF74713;
mem['h02E9] = 32'h06E12C23;
mem['h02EA] = 32'h00010613;
mem['h02EB] = 32'h0016C703;
mem['h02EC] = 32'h0026C583;
mem['h02ED] = 32'h00468693;
mem['h02EE] = 32'h00871713;
mem['h02EF] = 32'h01059593;
mem['h02F0] = 32'h00B74733;
mem['h02F1] = 32'hFFC6C583;
mem['h02F2] = 32'h00460613;
mem['h02F3] = 32'h00B74733;
mem['h02F4] = 32'hFFF6C583;
mem['h02F5] = 32'h01859593;
mem['h02F6] = 32'h00B74733;
mem['h02F7] = 32'hFEE62E23;
mem['h02F8] = 32'hFCDE16E3;
mem['h02F9] = 32'h04012903;
mem['h02FA] = 32'h05012603;
mem['h02FB] = 32'h06012A83;
mem['h02FC] = 32'h04412383;
mem['h02FD] = 32'h05412303;
mem['h02FE] = 32'h06412A03;
mem['h02FF] = 32'h04812983;
mem['h0300] = 32'h05812803;
mem['h0301] = 32'h07812703;
mem['h0302] = 32'h06812483;
mem['h0303] = 32'h04C12283;
mem['h0304] = 32'h05C12503;
mem['h0305] = 32'h07C12683;
mem['h0306] = 32'h06C12403;
mem['h0307] = 32'h08010F93;
mem['h0308] = 32'h000FC583;
mem['h0309] = 32'h010F8F93;
mem['h030A] = 32'h00259593;
mem['h030B] = 32'h12058593;
mem['h030C] = 32'h002585B3;
mem['h030D] = 32'hEE05AB03;
mem['h030E] = 32'h01660B33;
mem['h030F] = 32'h012B0B33;
mem['h0310] = 32'h011B45B3;
mem['h0311] = 32'h01059893;
mem['h0312] = 32'h0105D593;
mem['h0313] = 32'h0115E5B3;
mem['h0314] = 32'h01558AB3;
mem['h0315] = 32'h00CAC633;
mem['h0316] = 32'h00C65893;
mem['h0317] = 32'h01461613;
mem['h0318] = 32'h01166633;
mem['h0319] = 32'hFF1FC883;
mem['h031A] = 32'h00289893;
mem['h031B] = 32'h12088893;
mem['h031C] = 32'h002888B3;
mem['h031D] = 32'hEE08A903;
mem['h031E] = 32'h01260933;
mem['h031F] = 32'h01690933;
mem['h0320] = 32'h0125C5B3;
mem['h0321] = 32'h0085D893;
mem['h0322] = 32'h01859593;
mem['h0323] = 32'h0115E5B3;
mem['h0324] = 32'h00BA8AB3;
mem['h0325] = 32'h01564633;
mem['h0326] = 32'h00765893;
mem['h0327] = 32'h01961613;
mem['h0328] = 32'h01166633;
mem['h0329] = 32'hFF2FC883;
mem['h032A] = 32'h00289893;
mem['h032B] = 32'h12088893;
mem['h032C] = 32'h002888B3;
mem['h032D] = 32'hEE08A883;
mem['h032E] = 32'h011308B3;
mem['h032F] = 32'h007888B3;
mem['h0330] = 32'h00F8C7B3;
mem['h0331] = 32'h01079393;
mem['h0332] = 32'h0107D793;
mem['h0333] = 32'h0077E7B3;
mem['h0334] = 32'h01478A33;
mem['h0335] = 32'h006A4333;
mem['h0336] = 32'h00C35393;
mem['h0337] = 32'h01431313;
mem['h0338] = 32'h00736333;
mem['h0339] = 32'hFF3FC383;
mem['h033A] = 32'h00239393;
mem['h033B] = 32'h12038393;
mem['h033C] = 32'h002383B3;
mem['h033D] = 32'hEE03A383;
mem['h033E] = 32'h007303B3;
mem['h033F] = 32'h011383B3;
mem['h0340] = 32'h0077C7B3;
mem['h0341] = 32'h0087D893;
mem['h0342] = 32'h01879793;
mem['h0343] = 32'h0117E7B3;
mem['h0344] = 32'h00FA0A33;
mem['h0345] = 32'h01434333;
mem['h0346] = 32'h00735893;
mem['h0347] = 32'h01931313;
mem['h0348] = 32'h01136333;
mem['h0349] = 32'hFF4FC883;
mem['h034A] = 32'h00289893;
mem['h034B] = 32'h12088893;
mem['h034C] = 32'h002888B3;
mem['h034D] = 32'hEE08A883;
mem['h034E] = 32'h011808B3;
mem['h034F] = 32'h013888B3;
mem['h0350] = 32'h00E8C733;
mem['h0351] = 32'h01071993;
mem['h0352] = 32'h01075713;
mem['h0353] = 32'h01376733;
mem['h0354] = 32'h009704B3;
mem['h0355] = 32'h0104C833;
mem['h0356] = 32'h00C85993;
mem['h0357] = 32'h01481813;
mem['h0358] = 32'h01386833;
mem['h0359] = 32'hFF5FC983;
mem['h035A] = 32'h00299993;
mem['h035B] = 32'h12098993;
mem['h035C] = 32'h002989B3;
mem['h035D] = 32'hEE09A983;
mem['h035E] = 32'h013809B3;
mem['h035F] = 32'h011989B3;
mem['h0360] = 32'h01374733;
mem['h0361] = 32'h00875893;
mem['h0362] = 32'h01871713;
mem['h0363] = 32'h01176733;
mem['h0364] = 32'h00E484B3;
mem['h0365] = 32'h00984833;
mem['h0366] = 32'h00785893;
mem['h0367] = 32'h01981813;
mem['h0368] = 32'h01186833;
mem['h0369] = 32'hFF6FC883;
mem['h036A] = 32'h00289893;
mem['h036B] = 32'h12088893;
mem['h036C] = 32'h002888B3;
mem['h036D] = 32'hEE08A883;
mem['h036E] = 32'h011508B3;
mem['h036F] = 32'h005888B3;
mem['h0370] = 32'h00D8C6B3;
mem['h0371] = 32'h01069293;
mem['h0372] = 32'h0106D693;
mem['h0373] = 32'h0056E6B3;
mem['h0374] = 32'h00868433;
mem['h0375] = 32'h00A44533;
mem['h0376] = 32'h00C55293;
mem['h0377] = 32'h01451513;
mem['h0378] = 32'h00556533;
mem['h0379] = 32'hFF7FC283;
mem['h037A] = 32'h00229293;
mem['h037B] = 32'h12028293;
mem['h037C] = 32'h002282B3;
mem['h037D] = 32'hEE02A283;
mem['h037E] = 32'h005502B3;
mem['h037F] = 32'h011282B3;
mem['h0380] = 32'h0056C6B3;
mem['h0381] = 32'h0086D893;
mem['h0382] = 32'h01869693;
mem['h0383] = 32'h0116E6B3;
mem['h0384] = 32'h00D40433;
mem['h0385] = 32'h00854533;
mem['h0386] = 32'h00755893;
mem['h0387] = 32'h01951513;
mem['h0388] = 32'h01156533;
mem['h0389] = 32'hFF8FC883;
mem['h038A] = 32'h00289893;
mem['h038B] = 32'h12088893;
mem['h038C] = 32'h002888B3;
mem['h038D] = 32'hEE08A883;
mem['h038E] = 32'h01190933;
mem['h038F] = 32'h00690933;
mem['h0390] = 32'h0126C6B3;
mem['h0391] = 32'h01069893;
mem['h0392] = 32'h0106D693;
mem['h0393] = 32'h0116E6B3;
mem['h0394] = 32'h00D484B3;
mem['h0395] = 32'h00934333;
mem['h0396] = 32'h00C35893;
mem['h0397] = 32'h01431313;
mem['h0398] = 32'h01136333;
mem['h0399] = 32'hFF9FC883;
mem['h039A] = 32'h00289893;
mem['h039B] = 32'h12088893;
mem['h039C] = 32'h002888B3;
mem['h039D] = 32'hEE08A883;
mem['h039E] = 32'h01190933;
mem['h039F] = 32'h00690933;
mem['h03A0] = 32'h0126C6B3;
mem['h03A1] = 32'h0086D893;
mem['h03A2] = 32'h01869693;
mem['h03A3] = 32'h0116E6B3;
mem['h03A4] = 32'h00D484B3;
mem['h03A5] = 32'h00934333;
mem['h03A6] = 32'h00735893;
mem['h03A7] = 32'h01931313;
mem['h03A8] = 32'h01136333;
mem['h03A9] = 32'hFFAFC883;
mem['h03AA] = 32'h00289893;
mem['h03AB] = 32'h12088893;
mem['h03AC] = 32'h002888B3;
mem['h03AD] = 32'hEE08A883;
mem['h03AE] = 32'h011383B3;
mem['h03AF] = 32'h010383B3;
mem['h03B0] = 32'h0075C5B3;
mem['h03B1] = 32'h01059B13;
mem['h03B2] = 32'h0105D893;
mem['h03B3] = 32'h0168E8B3;
mem['h03B4] = 32'h01140433;
mem['h03B5] = 32'h00884833;
mem['h03B6] = 32'h00C85593;
mem['h03B7] = 32'h01481813;
mem['h03B8] = 32'h00B86833;
mem['h03B9] = 32'hFFBFC583;
mem['h03BA] = 32'h00259593;
mem['h03BB] = 32'h12058593;
mem['h03BC] = 32'h002585B3;
mem['h03BD] = 32'hEE05A583;
mem['h03BE] = 32'h00B383B3;
mem['h03BF] = 32'h010383B3;
mem['h03C0] = 32'h0078C8B3;
mem['h03C1] = 32'h0088D593;
mem['h03C2] = 32'h01889893;
mem['h03C3] = 32'h00B8E8B3;
mem['h03C4] = 32'h01140433;
mem['h03C5] = 32'h00884833;
mem['h03C6] = 32'h00785593;
mem['h03C7] = 32'h01981813;
mem['h03C8] = 32'h00B86833;
mem['h03C9] = 32'hFFCFC583;
mem['h03CA] = 32'h00259593;
mem['h03CB] = 32'h12058593;
mem['h03CC] = 32'h002585B3;
mem['h03CD] = 32'hEE05A583;
mem['h03CE] = 32'h00B989B3;
mem['h03CF] = 32'h00A989B3;
mem['h03D0] = 32'h0137C7B3;
mem['h03D1] = 32'h01079593;
mem['h03D2] = 32'h0107D793;
mem['h03D3] = 32'h00B7E7B3;
mem['h03D4] = 32'h00FA8AB3;
mem['h03D5] = 32'h01554533;
mem['h03D6] = 32'h00C55593;
mem['h03D7] = 32'h01451513;
mem['h03D8] = 32'h00B56533;
mem['h03D9] = 32'hFFDFC583;
mem['h03DA] = 32'h00259593;
mem['h03DB] = 32'h12058593;
mem['h03DC] = 32'h002585B3;
mem['h03DD] = 32'hEE05A583;
mem['h03DE] = 32'h00B989B3;
mem['h03DF] = 32'h00A989B3;
mem['h03E0] = 32'h0137C7B3;
mem['h03E1] = 32'h0087D593;
mem['h03E2] = 32'h01879793;
mem['h03E3] = 32'h00B7E7B3;
mem['h03E4] = 32'h00FA8AB3;
mem['h03E5] = 32'h01554533;
mem['h03E6] = 32'h00755593;
mem['h03E7] = 32'h01951513;
mem['h03E8] = 32'h00B56533;
mem['h03E9] = 32'hFFEFC583;
mem['h03EA] = 32'h00259593;
mem['h03EB] = 32'h12058593;
mem['h03EC] = 32'h002585B3;
mem['h03ED] = 32'hEE05A583;
mem['h03EE] = 32'h00B282B3;
mem['h03EF] = 32'h00C282B3;
mem['h03F0] = 32'h00574733;
mem['h03F1] = 32'h01071593;
mem['h03F2] = 32'h01075713;
mem['h03F3] = 32'h00B76733;
mem['h03F4] = 32'h00EA0A33;
mem['h03F5] = 32'h01464633;
mem['h03F6] = 32'h00C65593;
mem['h03F7] = 32'h01461613;
mem['h03F8] = 32'h00B66633;
mem['h03F9] = 32'hFFFFC583;
mem['h03FA] = 32'h00259593;
mem['h03FB] = 32'h12058593;
mem['h03FC] = 32'h002585B3;
mem['h03FD] = 32'hEE05A583;
mem['h03FE] = 32'h00B282B3;
mem['h03FF] = 32'h00C282B3;
mem['h0400] = 32'h00574733;
mem['h0401] = 32'h00875593;
mem['h0402] = 32'h01871713;
mem['h0403] = 32'h00B76733;
mem['h0404] = 32'h00EA0A33;
mem['h0405] = 32'h01464633;
mem['h0406] = 32'h00765593;
mem['h0407] = 32'h01961613;
mem['h0408] = 32'h00B66633;
mem['h0409] = 32'h12010593;
mem['h040A] = 32'hBFF59CE3;
mem['h040B] = 32'h05212023;
mem['h040C] = 32'h06D12E23;
mem['h040D] = 32'h06912423;
mem['h040E] = 32'h04612A23;
mem['h040F] = 32'h04712223;
mem['h0410] = 32'h07112823;
mem['h0411] = 32'h06812623;
mem['h0412] = 32'h05012C23;
mem['h0413] = 32'h05312423;
mem['h0414] = 32'h06F12A23;
mem['h0415] = 32'h07512023;
mem['h0416] = 32'h04A12E23;
mem['h0417] = 32'h04512623;
mem['h0418] = 32'h06E12C23;
mem['h0419] = 32'h07412223;
mem['h041A] = 32'h04C12823;
mem['h041B] = 32'h000E2783;
mem['h041C] = 32'h000EA703;
mem['h041D] = 32'h004E0E13;
mem['h041E] = 32'h004E8E93;
mem['h041F] = 32'h00E7C7B3;
mem['h0420] = 32'h01CEA703;
mem['h0421] = 32'h00E7C7B3;
mem['h0422] = 32'hFEFE2E23;
mem['h0423] = 32'hFFCF10E3;
mem['h0424] = 32'h13C12083;
mem['h0425] = 32'h13812403;
mem['h0426] = 32'h13412483;
mem['h0427] = 32'h13012903;
mem['h0428] = 32'h12C12983;
mem['h0429] = 32'h12812A03;
mem['h042A] = 32'h12412A83;
mem['h042B] = 32'h12012B03;
mem['h042C] = 32'h14010113;
mem['h042D] = 32'h00008067;
mem['h042E] = 32'h100096B7;
mem['h042F] = 32'hC246A703;
mem['h0430] = 32'h100017B7;
mem['h0431] = 32'hC2478793;
mem['h0432] = 32'h00F707B3;
mem['h0433] = 32'h00A70733;
mem['h0434] = 32'hC2E6A223;
mem['h0435] = 32'h000086B7;
mem['h0436] = 32'h00E6D463;
mem['h0437] = 32'h00100073;
mem['h0438] = 32'h00078513;
mem['h0439] = 32'h00008067;
mem['h043A] = 32'hFE010113;
mem['h043B] = 32'h00912A23;
mem['h043C] = 32'h00058493;
mem['h043D] = 32'h000055B7;
mem['h043E] = 32'h78458593;
mem['h043F] = 32'h00112E23;
mem['h0440] = 32'h00812C23;
mem['h0441] = 32'h01212823;
mem['h0442] = 32'h00050413;
mem['h0443] = 32'h8B8FF0EF;
mem['h0444] = 32'h00048593;
mem['h0445] = 32'h00040513;
mem['h0446] = 32'hFF1FE0EF;
mem['h0447] = 32'h02842783;
mem['h0448] = 32'h00249493;
mem['h0449] = 32'h000055B7;
mem['h044A] = 32'h009787B3;
mem['h044B] = 32'h0007A783;
mem['h044C] = 32'h00040513;
mem['h044D] = 32'h78858593;
mem['h044E] = 32'h0007A783;
mem['h044F] = 32'h0007A683;
mem['h0450] = 32'h0006D783;
mem['h0451] = 32'h00879713;
mem['h0452] = 32'h0087D793;
mem['h0453] = 32'h00F76733;
mem['h0454] = 32'h0006A783;
mem['h0455] = 32'h00E11723;
mem['h0456] = 32'h0187D693;
mem['h0457] = 32'h0107D793;
mem['h0458] = 32'h00D10623;
mem['h0459] = 32'h00F106A3;
mem['h045A] = 32'h85CFF0EF;
mem['h045B] = 32'h00C10593;
mem['h045C] = 32'h00040513;
mem['h045D] = 32'h894FF0EF;
mem['h045E] = 32'h02842783;
mem['h045F] = 32'h000055B7;
mem['h0460] = 32'h00040513;
mem['h0461] = 32'h009787B3;
mem['h0462] = 32'h0007A783;
mem['h0463] = 32'h79058593;
mem['h0464] = 32'h0047A783;
mem['h0465] = 32'h0007A683;
mem['h0466] = 32'h0006D783;
mem['h0467] = 32'h00879713;
mem['h0468] = 32'h0087D793;
mem['h0469] = 32'h00F76733;
mem['h046A] = 32'h0006A783;
mem['h046B] = 32'h00E11523;
mem['h046C] = 32'h0187D693;
mem['h046D] = 32'h0107D793;
mem['h046E] = 32'h00D10423;
mem['h046F] = 32'h00F104A3;
mem['h0470] = 32'h804FF0EF;
mem['h0471] = 32'h00810593;
mem['h0472] = 32'h00040513;
mem['h0473] = 32'h83CFF0EF;
mem['h0474] = 32'h02842783;
mem['h0475] = 32'h000055B7;
mem['h0476] = 32'h00040513;
mem['h0477] = 32'h009787B3;
mem['h0478] = 32'h0007A783;
mem['h0479] = 32'h79C58593;
mem['h047A] = 32'h0087A783;
mem['h047B] = 32'h0007A783;
mem['h047C] = 32'h0007A903;
mem['h047D] = 32'hFD1FE0EF;
mem['h047E] = 32'h00040513;
mem['h047F] = 32'h03F97913;
mem['h0480] = 32'h00090593;
mem['h0481] = 32'hF05FE0EF;
mem['h0482] = 32'h02842783;
mem['h0483] = 32'h000055B7;
mem['h0484] = 32'h00040513;
mem['h0485] = 32'h009787B3;
mem['h0486] = 32'h0007A783;
mem['h0487] = 32'h7AC58593;
mem['h0488] = 32'h00C7A783;
mem['h0489] = 32'h0007A783;
mem['h048A] = 32'h0007A483;
mem['h048B] = 32'hF99FE0EF;
mem['h048C] = 32'h00040513;
mem['h048D] = 32'h0074F493;
mem['h048E] = 32'h00048593;
mem['h048F] = 32'hECDFE0EF;
mem['h0490] = 32'h00040513;
mem['h0491] = 32'h01812403;
mem['h0492] = 32'h01C12083;
mem['h0493] = 32'h01412483;
mem['h0494] = 32'h01012903;
mem['h0495] = 32'h000065B7;
mem['h0496] = 32'hBF058593;
mem['h0497] = 32'h02010113;
mem['h0498] = 32'hF65FE06F;
mem['h0499] = 32'hFE010113;
mem['h049A] = 32'h00912A23;
mem['h049B] = 32'h00058493;
mem['h049C] = 32'h000055B7;
mem['h049D] = 32'h78458593;
mem['h049E] = 32'h00112E23;
mem['h049F] = 32'h00812C23;
mem['h04A0] = 32'h00050413;
mem['h04A1] = 32'hF41FE0EF;
mem['h04A2] = 32'h00048593;
mem['h04A3] = 32'h00040513;
mem['h04A4] = 32'hE79FE0EF;
mem['h04A5] = 32'h000055B7;
mem['h04A6] = 32'h00040513;
mem['h04A7] = 32'h7B458593;
mem['h04A8] = 32'hF25FE0EF;
mem['h04A9] = 32'h02C42783;
mem['h04AA] = 32'h00249493;
mem['h04AB] = 32'h00040513;
mem['h04AC] = 32'h009787B3;
mem['h04AD] = 32'h0007A783;
mem['h04AE] = 32'h00400613;
mem['h04AF] = 32'h0007A783;
mem['h04B0] = 32'h0007A783;
mem['h04B1] = 32'h0007D583;
mem['h04B2] = 32'hDD5FE0EF;
mem['h04B3] = 32'h02C42783;
mem['h04B4] = 32'h00800613;
mem['h04B5] = 32'h00040513;
mem['h04B6] = 32'h009787B3;
mem['h04B7] = 32'h0007A783;
mem['h04B8] = 32'h0047A783;
mem['h04B9] = 32'h0007A783;
mem['h04BA] = 32'h0007A583;
mem['h04BB] = 32'hDB1FE0EF;
mem['h04BC] = 32'h000055B7;
mem['h04BD] = 32'h00040513;
mem['h04BE] = 32'h7C458593;
mem['h04BF] = 32'hEC9FE0EF;
mem['h04C0] = 32'h02C42783;
mem['h04C1] = 32'h00C10593;
mem['h04C2] = 32'h00040513;
mem['h04C3] = 32'h009787B3;
mem['h04C4] = 32'h0007A783;
mem['h04C5] = 32'h0087A783;
mem['h04C6] = 32'h0007A683;
mem['h04C7] = 32'h0006D783;
mem['h04C8] = 32'h00879713;
mem['h04C9] = 32'h0087D793;
mem['h04CA] = 32'h00F76733;
mem['h04CB] = 32'h0006A783;
mem['h04CC] = 32'h00E11723;
mem['h04CD] = 32'h0187D693;
mem['h04CE] = 32'h0107D793;
mem['h04CF] = 32'h00D10623;
mem['h04D0] = 32'h00F106A3;
mem['h04D1] = 32'hEC5FE0EF;
mem['h04D2] = 32'h000055B7;
mem['h04D3] = 32'h00040513;
mem['h04D4] = 32'h7D458593;
mem['h04D5] = 32'hE71FE0EF;
mem['h04D6] = 32'h02C42783;
mem['h04D7] = 32'h00040513;
mem['h04D8] = 32'h009787B3;
mem['h04D9] = 32'h0007A783;
mem['h04DA] = 32'h00C7A783;
mem['h04DB] = 32'h0007A783;
mem['h04DC] = 32'h0007D583;
mem['h04DD] = 32'hD95FE0EF;
mem['h04DE] = 32'h000055B7;
mem['h04DF] = 32'h00040513;
mem['h04E0] = 32'h7E458593;
mem['h04E1] = 32'hE41FE0EF;
mem['h04E2] = 32'h02C42783;
mem['h04E3] = 32'h00800613;
mem['h04E4] = 32'h00040513;
mem['h04E5] = 32'h009787B3;
mem['h04E6] = 32'h0007A783;
mem['h04E7] = 32'h0107A783;
mem['h04E8] = 32'h0007A783;
mem['h04E9] = 32'h0007A583;
mem['h04EA] = 32'hCF5FE0EF;
mem['h04EB] = 32'h000055B7;
mem['h04EC] = 32'h00040513;
mem['h04ED] = 32'h7F458593;
mem['h04EE] = 32'hE0DFE0EF;
mem['h04EF] = 32'h02C42783;
mem['h04F0] = 32'h00040513;
mem['h04F1] = 32'h00400613;
mem['h04F2] = 32'h009787B3;
mem['h04F3] = 32'h0007A783;
mem['h04F4] = 32'h0147A783;
mem['h04F5] = 32'h0007A783;
mem['h04F6] = 32'h0007D583;
mem['h04F7] = 32'hCC1FE0EF;
mem['h04F8] = 32'h02C42783;
mem['h04F9] = 32'h00800613;
mem['h04FA] = 32'h00040513;
mem['h04FB] = 32'h009787B3;
mem['h04FC] = 32'h0007A783;
mem['h04FD] = 32'h0187A783;
mem['h04FE] = 32'h0007A783;
mem['h04FF] = 32'h0007A583;
mem['h0500] = 32'hC9DFE0EF;
mem['h0501] = 32'h000065B7;
mem['h0502] = 32'h00040513;
mem['h0503] = 32'h80858593;
mem['h0504] = 32'hDB5FE0EF;
mem['h0505] = 32'h02C42783;
mem['h0506] = 32'h00810593;
mem['h0507] = 32'h00040513;
mem['h0508] = 32'h009787B3;
mem['h0509] = 32'h0007A783;
mem['h050A] = 32'h01C7A783;
mem['h050B] = 32'h0007A683;
mem['h050C] = 32'h0006D783;
mem['h050D] = 32'h00879713;
mem['h050E] = 32'h0087D793;
mem['h050F] = 32'h00F76733;
mem['h0510] = 32'h0006A783;
mem['h0511] = 32'h00E11523;
mem['h0512] = 32'h0187D693;
mem['h0513] = 32'h0107D793;
mem['h0514] = 32'h00D10423;
mem['h0515] = 32'h00F104A3;
mem['h0516] = 32'hDB1FE0EF;
mem['h0517] = 32'h000065B7;
mem['h0518] = 32'h00040513;
mem['h0519] = 32'h81858593;
mem['h051A] = 32'hD5DFE0EF;
mem['h051B] = 32'h02C42783;
mem['h051C] = 32'h00040513;
mem['h051D] = 32'h009787B3;
mem['h051E] = 32'h0007A783;
mem['h051F] = 32'h0207A783;
mem['h0520] = 32'h0007A783;
mem['h0521] = 32'h0007D583;
mem['h0522] = 32'hC81FE0EF;
mem['h0523] = 32'h000065B7;
mem['h0524] = 32'h00040513;
mem['h0525] = 32'h82858593;
mem['h0526] = 32'hD2DFE0EF;
mem['h0527] = 32'h02C42783;
mem['h0528] = 32'h00800613;
mem['h0529] = 32'h00040513;
mem['h052A] = 32'h009787B3;
mem['h052B] = 32'h0007A783;
mem['h052C] = 32'h0247A783;
mem['h052D] = 32'h0007A783;
mem['h052E] = 32'h0007A583;
mem['h052F] = 32'hBE1FE0EF;
mem['h0530] = 32'h000065B7;
mem['h0531] = 32'h00040513;
mem['h0532] = 32'h83858593;
mem['h0533] = 32'hCF9FE0EF;
mem['h0534] = 32'h02C42783;
mem['h0535] = 32'h00040513;
mem['h0536] = 32'h00800613;
mem['h0537] = 32'h009787B3;
mem['h0538] = 32'h0007A783;
mem['h0539] = 32'h0287A783;
mem['h053A] = 32'h0007A783;
mem['h053B] = 32'h0007A583;
mem['h053C] = 32'hBADFE0EF;
mem['h053D] = 32'h02C42783;
mem['h053E] = 32'h00040513;
mem['h053F] = 32'h00800613;
mem['h0540] = 32'h009787B3;
mem['h0541] = 32'h0007A783;
mem['h0542] = 32'h02C7A783;
mem['h0543] = 32'h0007A783;
mem['h0544] = 32'h0007A583;
mem['h0545] = 32'hB89FE0EF;
mem['h0546] = 32'h02C42783;
mem['h0547] = 32'h00040513;
mem['h0548] = 32'h00800613;
mem['h0549] = 32'h009787B3;
mem['h054A] = 32'h0007A783;
mem['h054B] = 32'h0307A783;
mem['h054C] = 32'h0007A783;
mem['h054D] = 32'h0007A583;
mem['h054E] = 32'hB65FE0EF;
mem['h054F] = 32'h02C42783;
mem['h0550] = 32'h00040513;
mem['h0551] = 32'h00800613;
mem['h0552] = 32'h009787B3;
mem['h0553] = 32'h0007A783;
mem['h0554] = 32'h0347A783;
mem['h0555] = 32'h0007A783;
mem['h0556] = 32'h0007A583;
mem['h0557] = 32'hB41FE0EF;
mem['h0558] = 32'h02C42783;
mem['h0559] = 32'h00040513;
mem['h055A] = 32'h00800613;
mem['h055B] = 32'h009787B3;
mem['h055C] = 32'h0007A783;
mem['h055D] = 32'h0387A783;
mem['h055E] = 32'h0007A783;
mem['h055F] = 32'h0007A583;
mem['h0560] = 32'hB1DFE0EF;
mem['h0561] = 32'h02C42783;
mem['h0562] = 32'h00040513;
mem['h0563] = 32'h00800613;
mem['h0564] = 32'h009787B3;
mem['h0565] = 32'h0007A783;
mem['h0566] = 32'h03C7A783;
mem['h0567] = 32'h0007A783;
mem['h0568] = 32'h0007A583;
mem['h0569] = 32'hAF9FE0EF;
mem['h056A] = 32'h02C42783;
mem['h056B] = 32'h00040513;
mem['h056C] = 32'h00800613;
mem['h056D] = 32'h009787B3;
mem['h056E] = 32'h0007A783;
mem['h056F] = 32'h0407A783;
mem['h0570] = 32'h0007A783;
mem['h0571] = 32'h0007A583;
mem['h0572] = 32'hAD5FE0EF;
mem['h0573] = 32'h02C42783;
mem['h0574] = 32'h00800613;
mem['h0575] = 32'h00040513;
mem['h0576] = 32'h009787B3;
mem['h0577] = 32'h0007A783;
mem['h0578] = 32'h0447A783;
mem['h0579] = 32'h0007A783;
mem['h057A] = 32'h0007A583;
mem['h057B] = 32'hAB1FE0EF;
mem['h057C] = 32'h000065B7;
mem['h057D] = 32'h00040513;
mem['h057E] = 32'h85458593;
mem['h057F] = 32'hBC9FE0EF;
mem['h0580] = 32'h02C42783;
mem['h0581] = 32'h00040513;
mem['h0582] = 32'h00800613;
mem['h0583] = 32'h009787B3;
mem['h0584] = 32'h0007A783;
mem['h0585] = 32'h0487A783;
mem['h0586] = 32'h0007A783;
mem['h0587] = 32'h0007A583;
mem['h0588] = 32'hA7DFE0EF;
mem['h0589] = 32'h02C42783;
mem['h058A] = 32'h00040513;
mem['h058B] = 32'h00800613;
mem['h058C] = 32'h009787B3;
mem['h058D] = 32'h0007A783;
mem['h058E] = 32'h04C7A783;
mem['h058F] = 32'h0007A783;
mem['h0590] = 32'h0007A583;
mem['h0591] = 32'hA59FE0EF;
mem['h0592] = 32'h02C42783;
mem['h0593] = 32'h00040513;
mem['h0594] = 32'h00800613;
mem['h0595] = 32'h009787B3;
mem['h0596] = 32'h0007A783;
mem['h0597] = 32'h0507A783;
mem['h0598] = 32'h0007A783;
mem['h0599] = 32'h0007A583;
mem['h059A] = 32'hA35FE0EF;
mem['h059B] = 32'h02C42783;
mem['h059C] = 32'h00040513;
mem['h059D] = 32'h00800613;
mem['h059E] = 32'h009787B3;
mem['h059F] = 32'h0007A783;
mem['h05A0] = 32'h0547A783;
mem['h05A1] = 32'h0007A783;
mem['h05A2] = 32'h0007A583;
mem['h05A3] = 32'hA11FE0EF;
mem['h05A4] = 32'h02C42783;
mem['h05A5] = 32'h00040513;
mem['h05A6] = 32'h00800613;
mem['h05A7] = 32'h009787B3;
mem['h05A8] = 32'h0007A783;
mem['h05A9] = 32'h0587A783;
mem['h05AA] = 32'h0007A783;
mem['h05AB] = 32'h0007A583;
mem['h05AC] = 32'h9EDFE0EF;
mem['h05AD] = 32'h02C42783;
mem['h05AE] = 32'h00040513;
mem['h05AF] = 32'h00800613;
mem['h05B0] = 32'h009787B3;
mem['h05B1] = 32'h0007A783;
mem['h05B2] = 32'h05C7A783;
mem['h05B3] = 32'h0007A783;
mem['h05B4] = 32'h0007A583;
mem['h05B5] = 32'h9C9FE0EF;
mem['h05B6] = 32'h02C42783;
mem['h05B7] = 32'h00040513;
mem['h05B8] = 32'h00800613;
mem['h05B9] = 32'h009787B3;
mem['h05BA] = 32'h0007A783;
mem['h05BB] = 32'h0607A783;
mem['h05BC] = 32'h0007A783;
mem['h05BD] = 32'h0007A583;
mem['h05BE] = 32'h9A5FE0EF;
mem['h05BF] = 32'h02C42783;
mem['h05C0] = 32'h00800613;
mem['h05C1] = 32'h00040513;
mem['h05C2] = 32'h009787B3;
mem['h05C3] = 32'h0007A783;
mem['h05C4] = 32'h0647A783;
mem['h05C5] = 32'h0007A783;
mem['h05C6] = 32'h0007A583;
mem['h05C7] = 32'h981FE0EF;
mem['h05C8] = 32'h000065B7;
mem['h05C9] = 32'h00040513;
mem['h05CA] = 32'h87058593;
mem['h05CB] = 32'hA99FE0EF;
mem['h05CC] = 32'h02C42783;
mem['h05CD] = 32'h00040513;
mem['h05CE] = 32'h00800613;
mem['h05CF] = 32'h009787B3;
mem['h05D0] = 32'h0007A783;
mem['h05D1] = 32'h0687A783;
mem['h05D2] = 32'h0007A783;
mem['h05D3] = 32'h0007A583;
mem['h05D4] = 32'h94DFE0EF;
mem['h05D5] = 32'h02C42783;
mem['h05D6] = 32'h00800613;
mem['h05D7] = 32'h00040513;
mem['h05D8] = 32'h009787B3;
mem['h05D9] = 32'h0007A783;
mem['h05DA] = 32'h06C7A783;
mem['h05DB] = 32'h0007A783;
mem['h05DC] = 32'h0007A583;
mem['h05DD] = 32'h929FE0EF;
mem['h05DE] = 32'h000065B7;
mem['h05DF] = 32'h00040513;
mem['h05E0] = 32'h88858593;
mem['h05E1] = 32'hA41FE0EF;
mem['h05E2] = 32'h02C42783;
mem['h05E3] = 32'h00040513;
mem['h05E4] = 32'h00800613;
mem['h05E5] = 32'h009787B3;
mem['h05E6] = 32'h0007A783;
mem['h05E7] = 32'h0707A783;
mem['h05E8] = 32'h0007A783;
mem['h05E9] = 32'h0007A583;
mem['h05EA] = 32'h8F5FE0EF;
mem['h05EB] = 32'h02C42783;
mem['h05EC] = 32'h00040513;
mem['h05ED] = 32'h00800613;
mem['h05EE] = 32'h009787B3;
mem['h05EF] = 32'h0007A783;
mem['h05F0] = 32'h0747A783;
mem['h05F1] = 32'h0007A783;
mem['h05F2] = 32'h0007A583;
mem['h05F3] = 32'h8D1FE0EF;
mem['h05F4] = 32'h00040513;
mem['h05F5] = 32'h01812403;
mem['h05F6] = 32'h01C12083;
mem['h05F7] = 32'h01412483;
mem['h05F8] = 32'h000065B7;
mem['h05F9] = 32'hBF058593;
mem['h05FA] = 32'h02010113;
mem['h05FB] = 32'h9D9FE06F;
mem['h05FC] = 32'h000065B7;
mem['h05FD] = 32'hFF010113;
mem['h05FE] = 32'h8A058593;
mem['h05FF] = 32'h00112623;
mem['h0600] = 32'h00812423;
mem['h0601] = 32'h00912223;
mem['h0602] = 32'h00050413;
mem['h0603] = 32'h9B9FE0EF;
mem['h0604] = 32'h000065B7;
mem['h0605] = 32'h00040513;
mem['h0606] = 32'h8BC58593;
mem['h0607] = 32'h9A9FE0EF;
mem['h0608] = 32'h100005B7;
mem['h0609] = 32'h00058493;
mem['h060A] = 32'h00040513;
mem['h060B] = 32'h00058593;
mem['h060C] = 32'h9D9FE0EF;
mem['h060D] = 32'h000065B7;
mem['h060E] = 32'h00040513;
mem['h060F] = 32'h8D458593;
mem['h0610] = 32'h985FE0EF;
mem['h0611] = 32'h00448593;
mem['h0612] = 32'h00040513;
mem['h0613] = 32'h9BDFE0EF;
mem['h0614] = 32'h000065B7;
mem['h0615] = 32'h00040513;
mem['h0616] = 32'h8EC58593;
mem['h0617] = 32'h969FE0EF;
mem['h0618] = 32'h0084C583;
mem['h0619] = 32'h00200613;
mem['h061A] = 32'h00040513;
mem['h061B] = 32'h831FE0EF;
mem['h061C] = 32'h00040513;
mem['h061D] = 32'h03A00593;
mem['h061E] = 32'hFFCFE0EF;
mem['h061F] = 32'h0094C583;
mem['h0620] = 32'h00200613;
mem['h0621] = 32'h00040513;
mem['h0622] = 32'h815FE0EF;
mem['h0623] = 32'h00040513;
mem['h0624] = 32'h03A00593;
mem['h0625] = 32'hFE0FE0EF;
mem['h0626] = 32'h00A4C583;
mem['h0627] = 32'h00200613;
mem['h0628] = 32'h00040513;
mem['h0629] = 32'hFF8FE0EF;
mem['h062A] = 32'h00040513;
mem['h062B] = 32'h03A00593;
mem['h062C] = 32'hFC4FE0EF;
mem['h062D] = 32'h00B4C583;
mem['h062E] = 32'h00200613;
mem['h062F] = 32'h00040513;
mem['h0630] = 32'hFDCFE0EF;
mem['h0631] = 32'h00040513;
mem['h0632] = 32'h03A00593;
mem['h0633] = 32'hFA8FE0EF;
mem['h0634] = 32'h00C4C583;
mem['h0635] = 32'h00200613;
mem['h0636] = 32'h00040513;
mem['h0637] = 32'hFC0FE0EF;
mem['h0638] = 32'h00040513;
mem['h0639] = 32'h03A00593;
mem['h063A] = 32'hF8CFE0EF;
mem['h063B] = 32'h00D4C583;
mem['h063C] = 32'h00200613;
mem['h063D] = 32'h00040513;
mem['h063E] = 32'hFA4FE0EF;
mem['h063F] = 32'h000065B7;
mem['h0640] = 32'h00040513;
mem['h0641] = 32'h90458593;
mem['h0642] = 32'h8BDFE0EF;
mem['h0643] = 32'h00E48593;
mem['h0644] = 32'h00040513;
mem['h0645] = 32'h8F5FE0EF;
mem['h0646] = 32'h000065B7;
mem['h0647] = 32'h00040513;
mem['h0648] = 32'h91C58593;
mem['h0649] = 32'h8A1FE0EF;
mem['h064A] = 32'h0124C583;
mem['h064B] = 32'h00040513;
mem['h064C] = 32'hFD8FE0EF;
mem['h064D] = 32'h00040513;
mem['h064E] = 32'h00812403;
mem['h064F] = 32'h00C12083;
mem['h0650] = 32'h00412483;
mem['h0651] = 32'h000065B7;
mem['h0652] = 32'hBF058593;
mem['h0653] = 32'h01010113;
mem['h0654] = 32'h875FE06F;
mem['h0655] = 32'h00054783;
mem['h0656] = 32'h00A00713;
mem['h0657] = 32'h08E78063;
mem['h0658] = 32'h06078E63;
mem['h0659] = 32'h00000793;
mem['h065A] = 32'h00A00893;
mem['h065B] = 32'h00900313;
mem['h065C] = 32'h00500813;
mem['h065D] = 32'h00054703;
mem['h065E] = 32'h05171063;
mem['h065F] = 32'h04F67E63;
mem['h0660] = 32'h00008067;
mem['h0661] = 32'hFBF70693;
mem['h0662] = 32'h0FF6F693;
mem['h0663] = 32'h00D86A63;
mem['h0664] = 32'h00479793;
mem['h0665] = 32'hFC970713;
mem['h0666] = 32'h00F767B3;
mem['h0667] = 32'h0340006F;
mem['h0668] = 32'hF9F70693;
mem['h0669] = 32'h0FF6F693;
mem['h066A] = 32'h02D86A63;
mem['h066B] = 32'h00479793;
mem['h066C] = 32'hFA970713;
mem['h066D] = 32'hFE5FF06F;
mem['h066E] = 32'hFC0702E3;
mem['h066F] = 32'hFD070693;
mem['h0670] = 32'h0FF6FE13;
mem['h0671] = 32'hFDC360E3;
mem['h0672] = 32'h00479793;
mem['h0673] = 32'h00F6E7B3;
mem['h0674] = 32'h00150513;
mem['h0675] = 32'hFA1FF06F;
mem['h0676] = 32'h00F5A023;
mem['h0677] = 32'h00008067;
mem['h0678] = 32'h93010113;
mem['h0679] = 32'h6C812423;
mem['h067A] = 32'h6C112623;
mem['h067B] = 32'h6C912223;
mem['h067C] = 32'h6D212023;
mem['h067D] = 32'h6B312E23;
mem['h067E] = 32'h6B412C23;
mem['h067F] = 32'h6B512A23;
mem['h0680] = 32'h6B612823;
mem['h0681] = 32'h6B712623;
mem['h0682] = 32'h00050413;
mem['h0683] = 32'h00000793;
mem['h0684] = 32'h01F00713;
mem['h0685] = 32'h00F58533;
mem['h0686] = 32'h00054503;
mem['h0687] = 32'h00F106B3;
mem['h0688] = 32'h00178793;
mem['h0689] = 32'h00A68023;
mem['h068A] = 32'hFEE796E3;
mem['h068B] = 32'h01F5C783;
mem['h068C] = 32'h42010493;
mem['h068D] = 32'h02060593;
mem['h068E] = 32'h03F7F793;
mem['h068F] = 32'h0407E793;
mem['h0690] = 32'h00F10FA3;
mem['h0691] = 32'h00014783;
mem['h0692] = 32'h00048713;
mem['h0693] = 32'hFF87F793;
mem['h0694] = 32'h00F10023;
mem['h0695] = 32'h00164783;
mem['h0696] = 32'h00064683;
mem['h0697] = 32'h00260613;
mem['h0698] = 32'h00879793;
mem['h0699] = 32'h00D786B3;
mem['h069A] = 32'h00F6B7B3;
mem['h069B] = 32'h00D72023;
mem['h069C] = 32'h00F72223;
mem['h069D] = 32'h00870713;
mem['h069E] = 32'hFCB61EE3;
mem['h069F] = 32'h49812783;
mem['h06A0] = 32'h48012E23;
mem['h06A1] = 32'h08000713;
mem['h06A2] = 32'h01179793;
mem['h06A3] = 32'h0117D793;
mem['h06A4] = 32'h48F12C23;
mem['h06A5] = 32'h00000793;
mem['h06A6] = 32'h00F48633;
mem['h06A7] = 32'h00462583;
mem['h06A8] = 32'h00062503;
mem['h06A9] = 32'h0A010693;
mem['h06AA] = 32'h00F686B3;
mem['h06AB] = 32'h00B6A223;
mem['h06AC] = 32'h00A6A023;
mem['h06AD] = 32'h12010693;
mem['h06AE] = 32'h00F686B3;
mem['h06AF] = 32'h00000593;
mem['h06B0] = 32'h00000613;
mem['h06B1] = 32'h00B6A023;
mem['h06B2] = 32'h00C6A223;
mem['h06B3] = 32'h02010693;
mem['h06B4] = 32'h00F686B3;
mem['h06B5] = 32'h00B6A023;
mem['h06B6] = 32'h00C6A223;
mem['h06B7] = 32'h1A010693;
mem['h06B8] = 32'h00F686B3;
mem['h06B9] = 32'h00B6A023;
mem['h06BA] = 32'h00C6A223;
mem['h06BB] = 32'h00878793;
mem['h06BC] = 32'hFAE794E3;
mem['h06BD] = 32'h00100713;
mem['h06BE] = 32'h00000793;
mem['h06BF] = 32'h00006AB7;
mem['h06C0] = 32'h1AE12023;
mem['h06C1] = 32'h1AF12223;
mem['h06C2] = 32'h02E12023;
mem['h06C3] = 32'h02F12223;
mem['h06C4] = 32'h0FE00993;
mem['h06C5] = 32'h00000A13;
mem['h06C6] = 32'h6F0A8A93;
mem['h06C7] = 32'hFFF00B13;
mem['h06C8] = 32'h01DA1713;
mem['h06C9] = 32'h0039D793;
mem['h06CA] = 32'h00F767B3;
mem['h06CB] = 32'h6A078793;
mem['h06CC] = 32'h002787B3;
mem['h06CD] = 32'h9607C903;
mem['h06CE] = 32'h0079F793;
mem['h06CF] = 32'h0A010593;
mem['h06D0] = 32'h40F95933;
mem['h06D1] = 32'h00197913;
mem['h06D2] = 32'h00090613;
mem['h06D3] = 32'h02010513;
mem['h06D4] = 32'hCCDFE0EF;
mem['h06D5] = 32'h00090613;
mem['h06D6] = 32'h1A010593;
mem['h06D7] = 32'h12010513;
mem['h06D8] = 32'hCBDFE0EF;
mem['h06D9] = 32'h12010613;
mem['h06DA] = 32'h02010593;
mem['h06DB] = 32'h22010513;
mem['h06DC] = 32'hD71FE0EF;
mem['h06DD] = 32'h02010593;
mem['h06DE] = 32'h00058513;
mem['h06DF] = 32'h12010613;
mem['h06E0] = 32'hDA9FE0EF;
mem['h06E1] = 32'h1A010613;
mem['h06E2] = 32'h0A010593;
mem['h06E3] = 32'h12010513;
mem['h06E4] = 32'hD51FE0EF;
mem['h06E5] = 32'h0A010593;
mem['h06E6] = 32'h00058513;
mem['h06E7] = 32'h1A010613;
mem['h06E8] = 32'hD89FE0EF;
mem['h06E9] = 32'h22010613;
mem['h06EA] = 32'h00060593;
mem['h06EB] = 32'h1A010513;
mem['h06EC] = 32'hDC1FE0EF;
mem['h06ED] = 32'h02010613;
mem['h06EE] = 32'h00060593;
mem['h06EF] = 32'h2A010513;
mem['h06F0] = 32'hDB1FE0EF;
mem['h06F1] = 32'h02010613;
mem['h06F2] = 32'h00060513;
mem['h06F3] = 32'h12010593;
mem['h06F4] = 32'hDA1FE0EF;
mem['h06F5] = 32'h22010613;
mem['h06F6] = 32'h0A010593;
mem['h06F7] = 32'h12010513;
mem['h06F8] = 32'hD91FE0EF;
mem['h06F9] = 32'h12010613;
mem['h06FA] = 32'h02010593;
mem['h06FB] = 32'h22010513;
mem['h06FC] = 32'hCF1FE0EF;
mem['h06FD] = 32'h02010593;
mem['h06FE] = 32'h00058513;
mem['h06FF] = 32'h12010613;
mem['h0700] = 32'hD29FE0EF;
mem['h0701] = 32'h02010613;
mem['h0702] = 32'h00060593;
mem['h0703] = 32'h0A010513;
mem['h0704] = 32'hD61FE0EF;
mem['h0705] = 32'h2A010613;
mem['h0706] = 32'h1A010593;
mem['h0707] = 32'h12010513;
mem['h0708] = 32'hD09FE0EF;
mem['h0709] = 32'h000A8613;
mem['h070A] = 32'h12010593;
mem['h070B] = 32'h02010513;
mem['h070C] = 32'hD41FE0EF;
mem['h070D] = 32'h02010593;
mem['h070E] = 32'h00058513;
mem['h070F] = 32'h1A010613;
mem['h0710] = 32'hCA1FE0EF;
mem['h0711] = 32'h12010593;
mem['h0712] = 32'h00058513;
mem['h0713] = 32'h02010613;
mem['h0714] = 32'hD21FE0EF;
mem['h0715] = 32'h2A010613;
mem['h0716] = 32'h1A010593;
mem['h0717] = 32'h02010513;
mem['h0718] = 32'hD11FE0EF;
mem['h0719] = 32'h00048613;
mem['h071A] = 32'h0A010593;
mem['h071B] = 32'h1A010513;
mem['h071C] = 32'hD01FE0EF;
mem['h071D] = 32'h22010613;
mem['h071E] = 32'h00060593;
mem['h071F] = 32'h0A010513;
mem['h0720] = 32'hCF1FE0EF;
mem['h0721] = 32'h00090613;
mem['h0722] = 32'h0A010593;
mem['h0723] = 32'h02010513;
mem['h0724] = 32'hB8DFE0EF;
mem['h0725] = 32'h00090613;
mem['h0726] = 32'h1A010593;
mem['h0727] = 32'h12010513;
mem['h0728] = 32'hB7DFE0EF;
mem['h0729] = 32'h0019B793;
mem['h072A] = 32'hFFF98993;
mem['h072B] = 32'h40FA0A33;
mem['h072C] = 32'hE76998E3;
mem['h072D] = 32'hE73A16E3;
mem['h072E] = 32'h00048713;
mem['h072F] = 32'h00000793;
mem['h0730] = 32'h08000693;
mem['h0731] = 32'h02010613;
mem['h0732] = 32'h00F60633;
mem['h0733] = 32'h00062503;
mem['h0734] = 32'h00462583;
mem['h0735] = 32'h12010613;
mem['h0736] = 32'h00F60633;
mem['h0737] = 32'h08A72023;
mem['h0738] = 32'h08B72223;
mem['h0739] = 32'h00062503;
mem['h073A] = 32'h00462583;
mem['h073B] = 32'h0A010613;
mem['h073C] = 32'h00F60633;
mem['h073D] = 32'h10A72023;
mem['h073E] = 32'h10B72223;
mem['h073F] = 32'h00062503;
mem['h0740] = 32'h00462583;
mem['h0741] = 32'h1A010613;
mem['h0742] = 32'h00F60633;
mem['h0743] = 32'h18A72023;
mem['h0744] = 32'h18B72223;
mem['h0745] = 32'h00062503;
mem['h0746] = 32'h00462583;
mem['h0747] = 32'h00878793;
mem['h0748] = 32'h20A72023;
mem['h0749] = 32'h20B72223;
mem['h074A] = 32'h00870713;
mem['h074B] = 32'hF8D79CE3;
mem['h074C] = 32'h00048713;
mem['h074D] = 32'h00000793;
mem['h074E] = 32'h08000693;
mem['h074F] = 32'h10072503;
mem['h0750] = 32'h10472583;
mem['h0751] = 32'h3A010613;
mem['h0752] = 32'h00F60633;
mem['h0753] = 32'h00A62023;
mem['h0754] = 32'h00B62223;
mem['h0755] = 32'h00878793;
mem['h0756] = 32'h00870713;
mem['h0757] = 32'hFED790E3;
mem['h0758] = 32'h0FB00913;
mem['h0759] = 32'hFFD00993;
mem['h075A] = 32'h3A010613;
mem['h075B] = 32'h00060593;
mem['h075C] = 32'h00060513;
mem['h075D] = 32'hBFDFE0EF;
mem['h075E] = 32'hFFD97793;
mem['h075F] = 32'hFFF90913;
mem['h0760] = 32'hFE0784E3;
mem['h0761] = 32'h3A010593;
mem['h0762] = 32'h52010613;
mem['h0763] = 32'h00058513;
mem['h0764] = 32'hBE1FE0EF;
mem['h0765] = 32'hFD391AE3;
mem['h0766] = 32'h00048713;
mem['h0767] = 32'h00000793;
mem['h0768] = 32'h08000693;
mem['h0769] = 32'h3A010613;
mem['h076A] = 32'h00F60633;
mem['h076B] = 32'h00062503;
mem['h076C] = 32'h00462583;
mem['h076D] = 32'h00878793;
mem['h076E] = 32'h10A72023;
mem['h076F] = 32'h10B72223;
mem['h0770] = 32'h00870713;
mem['h0771] = 32'hFED790E3;
mem['h0772] = 32'h4A010593;
mem['h0773] = 32'h52010613;
mem['h0774] = 32'h00058513;
mem['h0775] = 32'hB9DFE0EF;
mem['h0776] = 32'h00000793;
mem['h0777] = 32'h08000713;
mem['h0778] = 32'h0804A503;
mem['h0779] = 32'h0844A583;
mem['h077A] = 32'h3A010693;
mem['h077B] = 32'h00F686B3;
mem['h077C] = 32'h00A6A023;
mem['h077D] = 32'h00B6A223;
mem['h077E] = 32'h00878793;
mem['h077F] = 32'h00848493;
mem['h0780] = 32'hFEE790E3;
mem['h0781] = 32'h3A010513;
mem['h0782] = 32'h8B5FE0EF;
mem['h0783] = 32'h3A010513;
mem['h0784] = 32'h8ADFE0EF;
mem['h0785] = 32'h3A010513;
mem['h0786] = 32'hFFFF09B7;
mem['h0787] = 32'hFFFF0A37;
mem['h0788] = 32'h000104B7;
mem['h0789] = 32'hFFFF8937;
mem['h078A] = 32'h895FE0EF;
mem['h078B] = 32'h00200A93;
mem['h078C] = 32'h01398993;
mem['h078D] = 32'h001A0A13;
mem['h078E] = 32'hFFF48493;
mem['h078F] = 32'h07800B93;
mem['h0790] = 32'h00190913;
mem['h0791] = 32'h00100B13;
mem['h0792] = 32'h3A012783;
mem['h0793] = 32'h3A412703;
mem['h0794] = 32'h00800513;
mem['h0795] = 32'h013786B3;
mem['h0796] = 32'h00F6B7B3;
mem['h0797] = 32'hFFF70713;
mem['h0798] = 32'h00E787B3;
mem['h0799] = 32'h32F12223;
mem['h079A] = 32'h32010793;
mem['h079B] = 32'h32D12023;
mem['h079C] = 32'h00078593;
mem['h079D] = 32'h3A010713;
mem['h079E] = 32'h00A706B3;
mem['h079F] = 32'h0006A703;
mem['h07A0] = 32'h0046A683;
mem['h07A1] = 32'h0007A803;
mem['h07A2] = 32'h01470633;
mem['h07A3] = 32'h00E63733;
mem['h07A4] = 32'hFFF68693;
mem['h07A5] = 32'h00D70733;
mem['h07A6] = 32'h01085693;
mem['h07A7] = 32'h0016F693;
mem['h07A8] = 32'h40D606B3;
mem['h07A9] = 32'h00D63633;
mem['h07AA] = 32'h40C70733;
mem['h07AB] = 32'h00987833;
mem['h07AC] = 32'h00D7A423;
mem['h07AD] = 32'h00E7A623;
mem['h07AE] = 32'h0107A023;
mem['h07AF] = 32'h0007A223;
mem['h07B0] = 32'h00850513;
mem['h07B1] = 32'h00878793;
mem['h07B2] = 32'hFB7516E3;
mem['h07B3] = 32'h41812783;
mem['h07B4] = 32'h41C12603;
mem['h07B5] = 32'h39012683;
mem['h07B6] = 32'h01278733;
mem['h07B7] = 32'h00F737B3;
mem['h07B8] = 32'hFFF60613;
mem['h07B9] = 32'h00C787B3;
mem['h07BA] = 32'h0106D613;
mem['h07BB] = 32'h00167613;
mem['h07BC] = 32'h40C70633;
mem['h07BD] = 32'h00C73733;
mem['h07BE] = 32'h40E787B3;
mem['h07BF] = 32'h38C12C23;
mem['h07C0] = 32'h38F12E23;
mem['h07C1] = 32'h01065613;
mem['h07C2] = 32'h01079793;
mem['h07C3] = 32'h00C7E633;
mem['h07C4] = 32'hFFF64613;
mem['h07C5] = 32'h0096F6B3;
mem['h07C6] = 32'h00167613;
mem['h07C7] = 32'h3A010513;
mem['h07C8] = 32'h38D12823;
mem['h07C9] = 32'h38012A23;
mem['h07CA] = 32'h8F5FE0EF;
mem['h07CB] = 32'h056A9A63;
mem['h07CC] = 32'h3A010793;
mem['h07CD] = 32'h02040693;
mem['h07CE] = 32'h0007A703;
mem['h07CF] = 32'h00240413;
mem['h07D0] = 32'h00878793;
mem['h07D1] = 32'hFEE40F23;
mem['h07D2] = 32'h00875713;
mem['h07D3] = 32'hFEE40FA3;
mem['h07D4] = 32'hFE8694E3;
mem['h07D5] = 32'h6CC12083;
mem['h07D6] = 32'h6C812403;
mem['h07D7] = 32'h6C412483;
mem['h07D8] = 32'h6C012903;
mem['h07D9] = 32'h6BC12983;
mem['h07DA] = 32'h6B812A03;
mem['h07DB] = 32'h6B412A83;
mem['h07DC] = 32'h6B012B03;
mem['h07DD] = 32'h6AC12B83;
mem['h07DE] = 32'h6D010113;
mem['h07DF] = 32'h00008067;
mem['h07E0] = 32'h00100A93;
mem['h07E1] = 32'hEC5FF06F;
mem['h07E2] = 32'hFF010113;
mem['h07E3] = 32'h00012623;
mem['h07E4] = 32'h00000793;
mem['h07E5] = 32'h00000713;
mem['h07E6] = 32'h00A00813;
mem['h07E7] = 32'h00900893;
mem['h07E8] = 32'h02E00313;
mem['h07E9] = 32'h00200E13;
mem['h07EA] = 32'h0FF00E93;
mem['h07EB] = 32'h00054683;
mem['h07EC] = 32'h05069863;
mem['h07ED] = 32'h00300693;
mem['h07EE] = 32'h06D71663;
mem['h07EF] = 32'h00C14703;
mem['h07F0] = 32'h00F581A3;
mem['h07F1] = 32'h00E58023;
mem['h07F2] = 32'h00D14703;
mem['h07F3] = 32'h00E580A3;
mem['h07F4] = 32'h00E14703;
mem['h07F5] = 32'h00E58123;
mem['h07F6] = 32'h04C0006F;
mem['h07F7] = 32'h04669463;
mem['h07F8] = 32'h04EE4263;
mem['h07F9] = 32'h01070693;
mem['h07FA] = 32'h002686B3;
mem['h07FB] = 32'hFEF68E23;
mem['h07FC] = 32'h00170713;
mem['h07FD] = 32'h00000793;
mem['h07FE] = 32'h00150513;
mem['h07FF] = 32'hFB1FF06F;
mem['h0800] = 32'hFA068AE3;
mem['h0801] = 32'hFD068613;
mem['h0802] = 32'h0FF67F13;
mem['h0803] = 32'hFDE8E8E3;
mem['h0804] = 32'h00279693;
mem['h0805] = 32'h00F687B3;
mem['h0806] = 32'h00179793;
mem['h0807] = 32'h00F607B3;
mem['h0808] = 32'hFCFEDCE3;
mem['h0809] = 32'h01010113;
mem['h080A] = 32'h00008067;
mem['h080B] = 32'h00052783;
mem['h080C] = 32'h0007A783;
mem['h080D] = 32'h0187A783;
mem['h080E] = 32'h0007A783;
mem['h080F] = 32'h0007A783;
mem['h0810] = 32'h0017F793;
mem['h0811] = 32'h1E078E63;
mem['h0812] = 32'h00052783;
mem['h0813] = 32'h0005C703;
mem['h0814] = 32'hFFFF8637;
mem['h0815] = 32'h0007A783;
mem['h0816] = 32'h00777713;
mem['h0817] = 32'hFFFF08B7;
mem['h0818] = 32'h0107A783;
mem['h0819] = 32'hFFF60613;
mem['h081A] = 32'h0007A683;
mem['h081B] = 32'h0006A783;
mem['h081C] = 32'hFF87F793;
mem['h081D] = 32'h00E7E7B3;
mem['h081E] = 32'h00F6A023;
mem['h081F] = 32'h00052783;
mem['h0820] = 32'h0015C703;
mem['h0821] = 32'h0007A783;
mem['h0822] = 32'h00777713;
mem['h0823] = 32'h00371713;
mem['h0824] = 32'h0107A783;
mem['h0825] = 32'h0007A683;
mem['h0826] = 32'h0006A783;
mem['h0827] = 32'hFC77F793;
mem['h0828] = 32'h00E7E7B3;
mem['h0829] = 32'h00F6A023;
mem['h082A] = 32'h00052783;
mem['h082B] = 32'h0025C703;
mem['h082C] = 32'h0007A783;
mem['h082D] = 32'h00177713;
mem['h082E] = 32'h00671713;
mem['h082F] = 32'h0107A783;
mem['h0830] = 32'h0007A683;
mem['h0831] = 32'h0006A783;
mem['h0832] = 32'hFBF7F793;
mem['h0833] = 32'h00E7E7B3;
mem['h0834] = 32'h00F6A023;
mem['h0835] = 32'h00052783;
mem['h0836] = 32'h0035C703;
mem['h0837] = 32'h0007A783;
mem['h0838] = 32'h00177713;
mem['h0839] = 32'h00771713;
mem['h083A] = 32'h0107A783;
mem['h083B] = 32'h0007A683;
mem['h083C] = 32'h0006A783;
mem['h083D] = 32'hF7F7F793;
mem['h083E] = 32'h00E7E7B3;
mem['h083F] = 32'h00F6A023;
mem['h0840] = 32'h00858713;
mem['h0841] = 32'h00000793;
mem['h0842] = 32'h00052683;
mem['h0843] = 32'h00072803;
mem['h0844] = 32'h01078793;
mem['h0845] = 32'h0006A683;
mem['h0846] = 32'h01070713;
mem['h0847] = 32'h0006A683;
mem['h0848] = 32'h0006A683;
mem['h0849] = 32'h0106A023;
mem['h084A] = 32'h00052683;
mem['h084B] = 32'hFF472803;
mem['h084C] = 32'h0006A683;
mem['h084D] = 32'h0046A683;
mem['h084E] = 32'h0006A683;
mem['h084F] = 32'h0106A023;
mem['h0850] = 32'h00052683;
mem['h0851] = 32'hFF872803;
mem['h0852] = 32'h0006A683;
mem['h0853] = 32'h0086A683;
mem['h0854] = 32'h0006A683;
mem['h0855] = 32'h0106A023;
mem['h0856] = 32'h00052683;
mem['h0857] = 32'hFFC72803;
mem['h0858] = 32'h0006A683;
mem['h0859] = 32'h00C6A683;
mem['h085A] = 32'h0006A683;
mem['h085B] = 32'h0106A023;
mem['h085C] = 32'h0045A683;
mem['h085D] = 32'h04D7FE63;
mem['h085E] = 32'h00052683;
mem['h085F] = 32'h0006A683;
mem['h0860] = 32'h0106A683;
mem['h0861] = 32'h0006A803;
mem['h0862] = 32'h00082683;
mem['h0863] = 32'h0116E6B3;
mem['h0864] = 32'h00D82023;
mem['h0865] = 32'h00052683;
mem['h0866] = 32'h0006A683;
mem['h0867] = 32'h0106A683;
mem['h0868] = 32'h0006A803;
mem['h0869] = 32'h00082683;
mem['h086A] = 32'h00C6F6B3;
mem['h086B] = 32'h00D82023;
mem['h086C] = 32'h00052683;
mem['h086D] = 32'h0006A683;
mem['h086E] = 32'h0146A683;
mem['h086F] = 32'h0006A803;
mem['h0870] = 32'h00082683;
mem['h0871] = 32'h0016E693;
mem['h0872] = 32'h00D82023;
mem['h0873] = 32'hF3DFF06F;
mem['h0874] = 32'h00052703;
mem['h0875] = 32'h40D787B3;
mem['h0876] = 32'h000106B7;
mem['h0877] = 32'h00072703;
mem['h0878] = 32'hFFF68693;
mem['h0879] = 32'h40F6D7B3;
mem['h087A] = 32'h01072703;
mem['h087B] = 32'h01079793;
mem['h087C] = 32'h00072603;
mem['h087D] = 32'h00062703;
mem['h087E] = 32'h00D77733;
mem['h087F] = 32'h00F767B3;
mem['h0880] = 32'h00F62023;
mem['h0881] = 32'h00052783;
mem['h0882] = 32'h000086B7;
mem['h0883] = 32'h0007A783;
mem['h0884] = 32'h0107A783;
mem['h0885] = 32'h0007A703;
mem['h0886] = 32'h00072783;
mem['h0887] = 32'h00D7E7B3;
mem['h0888] = 32'h00F72023;
mem['h0889] = 32'h00052783;
mem['h088A] = 32'h0007A783;
mem['h088B] = 32'h0147A783;
mem['h088C] = 32'h0007A703;
mem['h088D] = 32'h00072783;
mem['h088E] = 32'h0017E793;
mem['h088F] = 32'h00F72023;
mem['h0890] = 32'h00008067;
mem['h0891] = 32'hBB67B7B7;
mem['h0892] = 32'hF7010113;
mem['h0893] = 32'hE8578793;
mem['h0894] = 32'h04F12223;
mem['h0895] = 32'h3C6EF7B7;
mem['h0896] = 32'h37278793;
mem['h0897] = 32'h04F12423;
mem['h0898] = 32'hA54FF7B7;
mem['h0899] = 32'h53A78793;
mem['h089A] = 32'h04F12623;
mem['h089B] = 32'h510E57B7;
mem['h089C] = 32'h27F78793;
mem['h089D] = 32'h04F12823;
mem['h089E] = 32'h9B0577B7;
mem['h089F] = 32'h88C78793;
mem['h08A0] = 32'h04F12A23;
mem['h08A1] = 32'h1F83E7B7;
mem['h08A2] = 32'h9AB78793;
mem['h08A3] = 32'h04F12C23;
mem['h08A4] = 32'h5BE0D7B7;
mem['h08A5] = 32'hD1978793;
mem['h08A6] = 32'h04F12E23;
mem['h08A7] = 32'h6B08E7B7;
mem['h08A8] = 32'h64778793;
mem['h08A9] = 32'h04F12023;
mem['h08AA] = 32'h02000793;
mem['h08AB] = 32'h08812423;
mem['h08AC] = 32'h08912223;
mem['h08AD] = 32'h06F12623;
mem['h08AE] = 32'h08112623;
mem['h08AF] = 32'h09212023;
mem['h08B0] = 32'h07312E23;
mem['h08B1] = 32'h07412C23;
mem['h08B2] = 32'h00050493;
mem['h08B3] = 32'h00058413;
mem['h08B4] = 32'h06012023;
mem['h08B5] = 32'h06012223;
mem['h08B6] = 32'h06012423;
mem['h08B7] = 32'h00000793;
mem['h08B8] = 32'h04000713;
mem['h08B9] = 32'h00F106B3;
mem['h08BA] = 32'h00068023;
mem['h08BB] = 32'h00178793;
mem['h08BC] = 32'hFEE79AE3;
mem['h08BD] = 32'h00C40933;
mem['h08BE] = 32'h04000993;
mem['h08BF] = 32'h03F00A13;
mem['h08C0] = 32'h06812703;
mem['h08C1] = 32'h06012783;
mem['h08C2] = 32'h08891263;
mem['h08C3] = 32'h00F707B3;
mem['h08C4] = 32'h06F12023;
mem['h08C5] = 32'h00E7F863;
mem['h08C6] = 32'h06412783;
mem['h08C7] = 32'h00178793;
mem['h08C8] = 32'h06F12223;
mem['h08C9] = 32'h00070793;
mem['h08CA] = 32'h00000693;
mem['h08CB] = 32'h03F00613;
mem['h08CC] = 32'h0AF67663;
mem['h08CD] = 32'h02068063;
mem['h08CE] = 32'h04173693;
mem['h08CF] = 32'h00000793;
mem['h08D0] = 32'h00068663;
mem['h08D1] = 32'h04000793;
mem['h08D2] = 32'h40E787B3;
mem['h08D3] = 32'h00E787B3;
mem['h08D4] = 32'h06F12423;
mem['h08D5] = 32'h00100593;
mem['h08D6] = 32'h00010513;
mem['h08D7] = 32'hFA4FE0EF;
mem['h08D8] = 32'h06C12603;
mem['h08D9] = 32'h00000793;
mem['h08DA] = 32'h08C79463;
mem['h08DB] = 32'h08C12083;
mem['h08DC] = 32'h08812403;
mem['h08DD] = 32'h08412483;
mem['h08DE] = 32'h08012903;
mem['h08DF] = 32'h07C12983;
mem['h08E0] = 32'h07812A03;
mem['h08E1] = 32'h09010113;
mem['h08E2] = 32'h00008067;
mem['h08E3] = 32'h03371663;
mem['h08E4] = 32'h04078793;
mem['h08E5] = 32'h06F12023;
mem['h08E6] = 32'h00FA6863;
mem['h08E7] = 32'h06412783;
mem['h08E8] = 32'h00178793;
mem['h08E9] = 32'h06F12223;
mem['h08EA] = 32'h00000593;
mem['h08EB] = 32'h00010513;
mem['h08EC] = 32'hF50FE0EF;
mem['h08ED] = 32'h06012423;
mem['h08EE] = 32'h06812783;
mem['h08EF] = 32'h00140413;
mem['h08F0] = 32'h00178713;
mem['h08F1] = 32'h06E12423;
mem['h08F2] = 32'hFFF44703;
mem['h08F3] = 32'h07078793;
mem['h08F4] = 32'h002787B3;
mem['h08F5] = 32'hF8E78823;
mem['h08F6] = 32'hF29FF06F;
mem['h08F7] = 32'h00F106B3;
mem['h08F8] = 32'h00068023;
mem['h08F9] = 32'h00178793;
mem['h08FA] = 32'h00100693;
mem['h08FB] = 32'hF45FF06F;
mem['h08FC] = 32'hFFC7F713;
mem['h08FD] = 32'h07070713;
mem['h08FE] = 32'h00270733;
mem['h08FF] = 32'hFD072703;
mem['h0900] = 32'h0037F693;
mem['h0901] = 32'h00369693;
mem['h0902] = 32'h00F485B3;
mem['h0903] = 32'h00D75733;
mem['h0904] = 32'h00E58023;
mem['h0905] = 32'h00178793;
mem['h0906] = 32'hF51FF06F;
mem['h0907] = 32'h0FF5F593;
mem['h0908] = 32'h00000793;
mem['h0909] = 32'h00C79463;
mem['h090A] = 32'h00008067;
mem['h090B] = 32'h00F50733;
mem['h090C] = 32'h00B70023;
mem['h090D] = 32'h00178793;
mem['h090E] = 32'hFEDFF06F;
mem['h090F] = 32'h01452783;
mem['h0910] = 32'hFC010113;
mem['h0911] = 32'h02812C23;
mem['h0912] = 32'h02912A23;
mem['h0913] = 32'h02112E23;
mem['h0914] = 32'hC007F493;
mem['h0915] = 32'h01052683;
mem['h0916] = 32'h00050413;
mem['h0917] = 32'h02049263;
mem['h0918] = 32'h01852703;
mem['h0919] = 32'h01C52603;
mem['h091A] = 32'h00C76733;
mem['h091B] = 32'h00071A63;
mem['h091C] = 32'h02052703;
mem['h091D] = 32'h02452603;
mem['h091E] = 32'h00C76733;
mem['h091F] = 32'h06070263;
mem['h0920] = 32'h3FF7F793;
mem['h0921] = 32'h00000813;
mem['h0922] = 32'h00F42A23;
mem['h0923] = 32'h00000793;
mem['h0924] = 32'h00D42823;
mem['h0925] = 32'h00F42C23;
mem['h0926] = 32'h01042E23;
mem['h0927] = 32'h02F42023;
mem['h0928] = 32'h03042223;
mem['h0929] = 32'h02800613;
mem['h092A] = 32'h00000593;
mem['h092B] = 32'h00810513;
mem['h092C] = 32'hF6DFF0EF;
mem['h092D] = 32'h00500613;
mem['h092E] = 32'h00000693;
mem['h092F] = 32'h00000513;
mem['h0930] = 32'h0024D593;
mem['h0931] = 32'h16C030EF;
mem['h0932] = 32'h00A12423;
mem['h0933] = 32'h00B12623;
mem['h0934] = 32'h00810613;
mem['h0935] = 32'h00040593;
mem['h0936] = 32'h00040513;
mem['h0937] = 32'h934FE0EF;
mem['h0938] = 32'h01442783;
mem['h0939] = 32'h01042703;
mem['h093A] = 32'hFFF00693;
mem['h093B] = 32'h3FF7F793;
mem['h093C] = 32'h06D71263;
mem['h093D] = 32'h3FF00693;
mem['h093E] = 32'h04D79E63;
mem['h093F] = 32'h00842783;
mem['h0940] = 32'h04E79A63;
mem['h0941] = 32'h00C42703;
mem['h0942] = 32'h04F71663;
mem['h0943] = 32'h00442683;
mem['h0944] = 32'h00042783;
mem['h0945] = 32'h04E69063;
mem['h0946] = 32'hFFA00713;
mem['h0947] = 32'h02F77C63;
mem['h0948] = 32'h00578713;
mem['h0949] = 32'h00F737B3;
mem['h094A] = 32'hFFF78793;
mem['h094B] = 32'h00F42223;
mem['h094C] = 32'h00000793;
mem['h094D] = 32'h00E42023;
mem['h094E] = 32'h00000813;
mem['h094F] = 32'h00F42423;
mem['h0950] = 32'hFFF00713;
mem['h0951] = 32'h3FF00793;
mem['h0952] = 32'h01042623;
mem['h0953] = 32'h00E42823;
mem['h0954] = 32'h00F42A23;
mem['h0955] = 32'h03C12083;
mem['h0956] = 32'h03812403;
mem['h0957] = 32'h03412483;
mem['h0958] = 32'h04010113;
mem['h0959] = 32'h00008067;
mem['h095A] = 32'hFE010113;
mem['h095B] = 32'h01212823;
mem['h095C] = 32'h02800613;
mem['h095D] = 32'h00058913;
mem['h095E] = 32'h00000593;
mem['h095F] = 32'h00812C23;
mem['h0960] = 32'h01312623;
mem['h0961] = 32'h01412423;
mem['h0962] = 32'h00112E23;
mem['h0963] = 32'h00912A23;
mem['h0964] = 32'h00050993;
mem['h0965] = 32'h00000413;
mem['h0966] = 32'hE85FF0EF;
mem['h0967] = 32'h01000A13;
mem['h0968] = 32'h008907B3;
mem['h0969] = 32'h0007C503;
mem['h096A] = 32'h00747613;
mem['h096B] = 32'hFF847493;
mem['h096C] = 32'h00361613;
mem['h096D] = 32'h00000593;
mem['h096E] = 32'h01C030EF;
mem['h096F] = 32'h009984B3;
mem['h0970] = 32'h0004A783;
mem['h0971] = 32'h00140413;
mem['h0972] = 32'h00A7E733;
mem['h0973] = 32'h0044A783;
mem['h0974] = 32'h00E4A023;
mem['h0975] = 32'h00B7E7B3;
mem['h0976] = 32'h00F4A223;
mem['h0977] = 32'hFD4412E3;
mem['h0978] = 32'h01C12083;
mem['h0979] = 32'h01812403;
mem['h097A] = 32'h01412483;
mem['h097B] = 32'h01012903;
mem['h097C] = 32'h00C12983;
mem['h097D] = 32'h00812A03;
mem['h097E] = 32'h02010113;
mem['h097F] = 32'h00008067;
mem['h0980] = 32'h00000793;
mem['h0981] = 32'h00C79463;
mem['h0982] = 32'h00008067;
mem['h0983] = 32'h00F58733;
mem['h0984] = 32'h00074683;
mem['h0985] = 32'h00F50733;
mem['h0986] = 32'h00178793;
mem['h0987] = 32'h00D70023;
mem['h0988] = 32'hFE5FF06F;
mem['h0989] = 32'hF0010113;
mem['h098A] = 32'h0D712E23;
mem['h098B] = 32'h0D912A23;
mem['h098C] = 32'h0DA12823;
mem['h098D] = 32'h0DB12623;
mem['h098E] = 32'h61708BB7;
mem['h098F] = 32'h33206CB7;
mem['h0990] = 32'h79623D37;
mem['h0991] = 32'h6B206DB7;
mem['h0992] = 32'h0E912A23;
mem['h0993] = 32'h0F212823;
mem['h0994] = 32'h0F312623;
mem['h0995] = 32'h0F412423;
mem['h0996] = 32'h0F512223;
mem['h0997] = 32'h0F612023;
mem['h0998] = 32'h0E112E23;
mem['h0999] = 32'h0E812C23;
mem['h099A] = 32'h0D812C23;
mem['h099B] = 32'h00050913;
mem['h099C] = 32'h00058993;
mem['h099D] = 32'h00060493;
mem['h099E] = 32'h00068B13;
mem['h099F] = 32'h00070A13;
mem['h09A0] = 32'h00078A93;
mem['h09A1] = 32'h865B8B93;
mem['h09A2] = 32'h46EC8C93;
mem['h09A3] = 32'hD32D0D13;
mem['h09A4] = 32'h574D8D93;
mem['h09A5] = 32'h04049063;
mem['h09A6] = 32'h0FC12083;
mem['h09A7] = 32'h0F812403;
mem['h09A8] = 32'h0F412483;
mem['h09A9] = 32'h0F012903;
mem['h09AA] = 32'h0EC12983;
mem['h09AB] = 32'h0E812A03;
mem['h09AC] = 32'h0E412A83;
mem['h09AD] = 32'h0E012B03;
mem['h09AE] = 32'h0DC12B83;
mem['h09AF] = 32'h0D812C03;
mem['h09B0] = 32'h0D412C83;
mem['h09B1] = 32'h0D012D03;
mem['h09B2] = 32'h0CC12D83;
mem['h09B3] = 32'h10010113;
mem['h09B4] = 32'h00008067;
mem['h09B5] = 32'h04010713;
mem['h09B6] = 32'h05712023;
mem['h09B7] = 32'h05912223;
mem['h09B8] = 32'h05A12423;
mem['h09B9] = 32'h05B12623;
mem['h09BA] = 32'h00000793;
mem['h09BB] = 32'h00070C13;
mem['h09BC] = 32'h02000693;
mem['h09BD] = 32'h00FB0633;
mem['h09BE] = 32'h00062603;
mem['h09BF] = 32'h00478793;
mem['h09C0] = 32'h00470713;
mem['h09C1] = 32'h00C72623;
mem['h09C2] = 32'hFED796E3;
mem['h09C3] = 32'h000A2783;
mem['h09C4] = 32'h04000613;
mem['h09C5] = 32'h000C0593;
mem['h09C6] = 32'h06F12A23;
mem['h09C7] = 32'h004A2783;
mem['h09C8] = 32'h08010513;
mem['h09C9] = 32'h07512823;
mem['h09CA] = 32'h06F12C23;
mem['h09CB] = 32'h008A2783;
mem['h09CC] = 32'h00A00413;
mem['h09CD] = 32'h06F12E23;
mem['h09CE] = 32'hEC9FF0EF;
mem['h09CF] = 32'h0B010693;
mem['h09D0] = 32'h0A010613;
mem['h09D1] = 32'h09010593;
mem['h09D2] = 32'h08010513;
mem['h09D3] = 32'hE2DFD0EF;
mem['h09D4] = 32'h0B410693;
mem['h09D5] = 32'h0A410613;
mem['h09D6] = 32'h09410593;
mem['h09D7] = 32'h08410513;
mem['h09D8] = 32'hE19FD0EF;
mem['h09D9] = 32'h0B810693;
mem['h09DA] = 32'h0A810613;
mem['h09DB] = 32'h09810593;
mem['h09DC] = 32'h08810513;
mem['h09DD] = 32'hE05FD0EF;
mem['h09DE] = 32'h0BC10693;
mem['h09DF] = 32'h0AC10613;
mem['h09E0] = 32'h09C10593;
mem['h09E1] = 32'h08C10513;
mem['h09E2] = 32'hDF1FD0EF;
mem['h09E3] = 32'h0BC10693;
mem['h09E4] = 32'h0A810613;
mem['h09E5] = 32'h09410593;
mem['h09E6] = 32'h08010513;
mem['h09E7] = 32'hDDDFD0EF;
mem['h09E8] = 32'h0B010693;
mem['h09E9] = 32'h0AC10613;
mem['h09EA] = 32'h09810593;
mem['h09EB] = 32'h08410513;
mem['h09EC] = 32'hDC9FD0EF;
mem['h09ED] = 32'h0B410693;
mem['h09EE] = 32'h0A010613;
mem['h09EF] = 32'h09C10593;
mem['h09F0] = 32'h08810513;
mem['h09F1] = 32'hDB5FD0EF;
mem['h09F2] = 32'h0B810693;
mem['h09F3] = 32'h0A410613;
mem['h09F4] = 32'h09010593;
mem['h09F5] = 32'h08C10513;
mem['h09F6] = 32'hFFF40413;
mem['h09F7] = 32'hD9DFD0EF;
mem['h09F8] = 32'hF4041EE3;
mem['h09F9] = 32'h00000613;
mem['h09FA] = 32'h04000713;
mem['h09FB] = 32'h08010793;
mem['h09FC] = 32'h00C787B3;
mem['h09FD] = 32'h00CC05B3;
mem['h09FE] = 32'h0007A783;
mem['h09FF] = 32'h0005A583;
mem['h0A00] = 32'h00C106B3;
mem['h0A01] = 32'h00460613;
mem['h0A02] = 32'h00B787B3;
mem['h0A03] = 32'h00F6A023;
mem['h0A04] = 32'hFCE61EE3;
mem['h0A05] = 32'h00048793;
mem['h0A06] = 32'h00967463;
mem['h0A07] = 32'h04000793;
mem['h0A08] = 32'h00898733;
mem['h0A09] = 32'h00810633;
mem['h0A0A] = 32'h00074703;
mem['h0A0B] = 32'h00064603;
mem['h0A0C] = 32'h008906B3;
mem['h0A0D] = 32'h00140413;
mem['h0A0E] = 32'h00C74733;
mem['h0A0F] = 32'h00E68023;
mem['h0A10] = 32'hFE8790E3;
mem['h0A11] = 32'h001A8A93;
mem['h0A12] = 32'h40F484B3;
mem['h0A13] = 32'h00F90933;
mem['h0A14] = 32'h00F989B3;
mem['h0A15] = 32'hE41FF06F;
mem['h0A16] = 32'hF8010113;
mem['h0A17] = 32'h07412423;
mem['h0A18] = 32'h07512223;
mem['h0A19] = 32'h00A12623;
mem['h0A1A] = 32'h00058A13;
mem['h0A1B] = 32'h00060A93;
mem['h0A1C] = 32'h00000593;
mem['h0A1D] = 32'h02800613;
mem['h0A1E] = 32'h01810513;
mem['h0A1F] = 32'h05812C23;
mem['h0A20] = 32'h05A12823;
mem['h0A21] = 32'h05B12623;
mem['h0A22] = 32'h06112E23;
mem['h0A23] = 32'h06812C23;
mem['h0A24] = 32'h06912A23;
mem['h0A25] = 32'h07212823;
mem['h0A26] = 32'h07312623;
mem['h0A27] = 32'h07612023;
mem['h0A28] = 32'h05712E23;
mem['h0A29] = 32'h05912A23;
mem['h0A2A] = 32'h01810D13;
mem['h0A2B] = 32'hB71FF0EF;
mem['h0A2C] = 32'h00000C13;
mem['h0A2D] = 32'h00500D93;
mem['h0A2E] = 32'h003C1793;
mem['h0A2F] = 32'h00FA07B3;
mem['h0A30] = 32'h0007A903;
mem['h0A31] = 32'h0047A983;
mem['h0A32] = 32'h000D0B93;
mem['h0A33] = 32'h00000C93;
mem['h0A34] = 32'h00000413;
mem['h0A35] = 32'h00000B13;
mem['h0A36] = 32'h418D84B3;
mem['h0A37] = 32'h003C9793;
mem['h0A38] = 32'h00FA87B3;
mem['h0A39] = 32'h0007A603;
mem['h0A3A] = 32'h0047A683;
mem['h0A3B] = 32'h00090513;
mem['h0A3C] = 32'h00098593;
mem['h0A3D] = 32'h53D020EF;
mem['h0A3E] = 32'h000BA703;
mem['h0A3F] = 32'h004BA683;
mem['h0A40] = 32'h00058893;
mem['h0A41] = 32'h00A70733;
mem['h0A42] = 32'h00B686B3;
mem['h0A43] = 32'h00A737B3;
mem['h0A44] = 32'h00D787B3;
mem['h0A45] = 32'h00870633;
mem['h0A46] = 32'h016785B3;
mem['h0A47] = 32'h00E636B3;
mem['h0A48] = 32'h00B686B3;
mem['h0A49] = 32'h00050313;
mem['h0A4A] = 32'h00100593;
mem['h0A4B] = 32'h0166E863;
mem['h0A4C] = 32'h00DB1463;
mem['h0A4D] = 32'h00866463;
mem['h0A4E] = 32'h00000593;
mem['h0A4F] = 32'h00100413;
mem['h0A50] = 32'h0117E863;
mem['h0A51] = 32'h00F89463;
mem['h0A52] = 32'h00676463;
mem['h0A53] = 32'h00000413;
mem['h0A54] = 32'h00858433;
mem['h0A55] = 32'h00CBA023;
mem['h0A56] = 32'h00DBA223;
mem['h0A57] = 32'h001C8C93;
mem['h0A58] = 32'h00B43B33;
mem['h0A59] = 32'h008B8B93;
mem['h0A5A] = 32'hF7949AE3;
mem['h0A5B] = 32'h001C0C13;
mem['h0A5C] = 32'h008D0D13;
mem['h0A5D] = 32'hF5BC12E3;
mem['h0A5E] = 32'h00C12503;
mem['h0A5F] = 32'h01810593;
mem['h0A60] = 32'h02800613;
mem['h0A61] = 32'hC7DFF0EF;
mem['h0A62] = 32'h07C12083;
mem['h0A63] = 32'h07812403;
mem['h0A64] = 32'h07412483;
mem['h0A65] = 32'h07012903;
mem['h0A66] = 32'h06C12983;
mem['h0A67] = 32'h06812A03;
mem['h0A68] = 32'h06412A83;
mem['h0A69] = 32'h06012B03;
mem['h0A6A] = 32'h05C12B83;
mem['h0A6B] = 32'h05812C03;
mem['h0A6C] = 32'h05412C83;
mem['h0A6D] = 32'h05012D03;
mem['h0A6E] = 32'h04C12D83;
mem['h0A6F] = 32'h08010113;
mem['h0A70] = 32'h00008067;
mem['h0A71] = 32'hEE010113;
mem['h0A72] = 32'h11212823;
mem['h0A73] = 32'h11412423;
mem['h0A74] = 32'h00060913;
mem['h0A75] = 32'h00050A13;
mem['h0A76] = 32'h01000613;
mem['h0A77] = 32'h01810513;
mem['h0A78] = 32'h10112E23;
mem['h0A79] = 32'h10812C23;
mem['h0A7A] = 32'h10912A23;
mem['h0A7B] = 32'h00068413;
mem['h0A7C] = 32'h00058493;
mem['h0A7D] = 32'h11312623;
mem['h0A7E] = 32'h11512223;
mem['h0A7F] = 32'hC05FF0EF;
mem['h0A80] = 32'h01048593;
mem['h0A81] = 32'h01000613;
mem['h0A82] = 32'h00810513;
mem['h0A83] = 32'hBF5FF0EF;
mem['h0A84] = 32'h01B14783;
mem['h0A85] = 32'h02800613;
mem['h0A86] = 32'h00000593;
mem['h0A87] = 32'h00F7F793;
mem['h0A88] = 32'h00F10DA3;
mem['h0A89] = 32'h01F14783;
mem['h0A8A] = 32'h03810513;
mem['h0A8B] = 32'h00445A93;
mem['h0A8C] = 32'h00F7F793;
mem['h0A8D] = 32'h00F10FA3;
mem['h0A8E] = 32'h02314783;
mem['h0A8F] = 32'h00F47493;
mem['h0A90] = 32'h00000993;
mem['h0A91] = 32'h00F7F793;
mem['h0A92] = 32'h02F101A3;
mem['h0A93] = 32'h02714783;
mem['h0A94] = 32'h00F7F793;
mem['h0A95] = 32'h02F103A3;
mem['h0A96] = 32'h01C14783;
mem['h0A97] = 32'hFFC7F793;
mem['h0A98] = 32'h00F10E23;
mem['h0A99] = 32'h02014783;
mem['h0A9A] = 32'hFFC7F793;
mem['h0A9B] = 32'h02F10023;
mem['h0A9C] = 32'h02414783;
mem['h0A9D] = 32'hFFC7F793;
mem['h0A9E] = 32'h02F10223;
mem['h0A9F] = 32'h9A1FF0EF;
mem['h0AA0] = 32'h01810593;
mem['h0AA1] = 32'h08810513;
mem['h0AA2] = 32'hAE1FF0EF;
mem['h0AA3] = 32'h00810593;
mem['h0AA4] = 32'h06010513;
mem['h0AA5] = 32'hAD5FF0EF;
mem['h0AA6] = 32'h0D599263;
mem['h0AA7] = 32'h06048E63;
mem['h0AA8] = 32'hFF047593;
mem['h0AA9] = 32'h00048613;
mem['h0AAA] = 32'h00B905B3;
mem['h0AAB] = 32'h02810513;
mem['h0AAC] = 32'h02012423;
mem['h0AAD] = 32'h02012623;
mem['h0AAE] = 32'h02012823;
mem['h0AAF] = 32'h02012A23;
mem['h0AB0] = 32'hB41FF0EF;
mem['h0AB1] = 32'h10048793;
mem['h0AB2] = 32'h002784B3;
mem['h0AB3] = 32'h02810593;
mem['h0AB4] = 32'h00100793;
mem['h0AB5] = 32'h0D810513;
mem['h0AB6] = 32'hF2F48423;
mem['h0AB7] = 32'hA8DFF0EF;
mem['h0AB8] = 32'h03810593;
mem['h0AB9] = 32'h00058513;
mem['h0ABA] = 32'h0D810613;
mem['h0ABB] = 32'hB25FD0EF;
mem['h0ABC] = 32'h02800613;
mem['h0ABD] = 32'h03810593;
mem['h0ABE] = 32'h0B010513;
mem['h0ABF] = 32'hB05FF0EF;
mem['h0AC0] = 32'h03810513;
mem['h0AC1] = 32'h08810613;
mem['h0AC2] = 32'h0B010593;
mem['h0AC3] = 32'hD4DFF0EF;
mem['h0AC4] = 32'h03810513;
mem['h0AC5] = 32'h929FF0EF;
mem['h0AC6] = 32'h03810593;
mem['h0AC7] = 32'h06010613;
mem['h0AC8] = 32'h00058513;
mem['h0AC9] = 32'hAEDFD0EF;
mem['h0ACA] = 32'h03810593;
mem['h0ACB] = 32'h000A0513;
mem['h0ACC] = 32'h01000613;
mem['h0ACD] = 32'hACDFF0EF;
mem['h0ACE] = 32'h11C12083;
mem['h0ACF] = 32'h11812403;
mem['h0AD0] = 32'h11412483;
mem['h0AD1] = 32'h11012903;
mem['h0AD2] = 32'h10C12983;
mem['h0AD3] = 32'h10812A03;
mem['h0AD4] = 32'h10412A83;
mem['h0AD5] = 32'h12010113;
mem['h0AD6] = 32'h00008067;
mem['h0AD7] = 32'h00499593;
mem['h0AD8] = 32'h00B905B3;
mem['h0AD9] = 32'h0D810513;
mem['h0ADA] = 32'hA01FF0EF;
mem['h0ADB] = 32'h0E812783;
mem['h0ADC] = 32'h03810593;
mem['h0ADD] = 32'h00058513;
mem['h0ADE] = 32'h0017E793;
mem['h0ADF] = 32'h0D810613;
mem['h0AE0] = 32'h0EF12423;
mem['h0AE1] = 32'hA8DFD0EF;
mem['h0AE2] = 32'h02800613;
mem['h0AE3] = 32'h03810593;
mem['h0AE4] = 32'h0B010513;
mem['h0AE5] = 32'hA6DFF0EF;
mem['h0AE6] = 32'h08810613;
mem['h0AE7] = 32'h0B010593;
mem['h0AE8] = 32'h03810513;
mem['h0AE9] = 32'hCB5FF0EF;
mem['h0AEA] = 32'h03810513;
mem['h0AEB] = 32'h891FF0EF;
mem['h0AEC] = 32'h00198993;
mem['h0AED] = 32'hEE5FF06F;
mem['h0AEE] = 32'hFA010113;
mem['h0AEF] = 32'h04812C23;
mem['h0AF0] = 32'h00B12623;
mem['h0AF1] = 32'h00050413;
mem['h0AF2] = 32'h00C12423;
mem['h0AF3] = 32'h00000593;
mem['h0AF4] = 32'h04000613;
mem['h0AF5] = 32'h01010513;
mem['h0AF6] = 32'h04112E23;
mem['h0AF7] = 32'h841FF0EF;
mem['h0AF8] = 32'h00812703;
mem['h0AF9] = 32'h00C12683;
mem['h0AFA] = 32'h01010593;
mem['h0AFB] = 32'h00058513;
mem['h0AFC] = 32'h00000793;
mem['h0AFD] = 32'h04000613;
mem['h0AFE] = 32'hA2DFF0EF;
mem['h0AFF] = 32'h01010593;
mem['h0B00] = 32'h00040513;
mem['h0B01] = 32'h02000613;
mem['h0B02] = 32'h9F9FF0EF;
mem['h0B03] = 32'h05C12083;
mem['h0B04] = 32'h05812403;
mem['h0B05] = 32'h06010113;
mem['h0B06] = 32'h00008067;
mem['h0B07] = 32'hF5010113;
mem['h0B08] = 32'h0A812423;
mem['h0B09] = 32'h0B212023;
mem['h0B0A] = 32'h09312E23;
mem['h0B0B] = 32'h00C10413;
mem['h0B0C] = 32'h6C0799B7;
mem['h0B0D] = 32'h5D589937;
mem['h0B0E] = 32'h0A912223;
mem['h0B0F] = 32'h09412C23;
mem['h0B10] = 32'h09512A23;
mem['h0B11] = 32'h09612823;
mem['h0B12] = 32'h0A112623;
mem['h0B13] = 32'h00050493;
mem['h0B14] = 32'h04C10A93;
mem['h0B15] = 32'h00040A13;
mem['h0B16] = 32'h96598993;
mem['h0B17] = 32'hB6590913;
mem['h0B18] = 32'h3E700B13;
mem['h0B19] = 32'hC00027F3;
mem['h0B1A] = 32'h0077D513;
mem['h0B1B] = 32'h00F54533;
mem['h0B1C] = 32'h00098593;
mem['h0B1D] = 32'h199020EF;
mem['h0B1E] = 32'h00B55793;
mem['h0B1F] = 32'h00A7C7B3;
mem['h0B20] = 32'h012787B3;
mem['h0B21] = 32'h00F42023;
mem['h0B22] = 32'h00012423;
mem['h0B23] = 32'h00812783;
mem['h0B24] = 32'h08FB5663;
mem['h0B25] = 32'h00440413;
mem['h0B26] = 32'hFD5416E3;
mem['h0B27] = 32'h00410913;
mem['h0B28] = 32'h000A0593;
mem['h0B29] = 32'h04000613;
mem['h0B2A] = 32'h00040513;
mem['h0B2B] = 32'h01212223;
mem['h0B2C] = 32'h951FF0EF;
mem['h0B2D] = 32'h00090593;
mem['h0B2E] = 32'h00400613;
mem['h0B2F] = 32'h08C10513;
mem['h0B30] = 32'h941FF0EF;
mem['h0B31] = 32'h00040593;
mem['h0B32] = 32'h00048513;
mem['h0B33] = 32'h04400613;
mem['h0B34] = 32'hD74FF0EF;
mem['h0B35] = 32'h04000613;
mem['h0B36] = 32'h00000593;
mem['h0B37] = 32'h000A0513;
mem['h0B38] = 32'hF3CFF0EF;
mem['h0B39] = 32'h00040513;
mem['h0B3A] = 32'h04400613;
mem['h0B3B] = 32'h00000593;
mem['h0B3C] = 32'hF2CFF0EF;
mem['h0B3D] = 32'h0AC12083;
mem['h0B3E] = 32'h0A812403;
mem['h0B3F] = 32'h0A412483;
mem['h0B40] = 32'h0A012903;
mem['h0B41] = 32'h09C12983;
mem['h0B42] = 32'h09812A03;
mem['h0B43] = 32'h09412A83;
mem['h0B44] = 32'h09012B03;
mem['h0B45] = 32'h0B010113;
mem['h0B46] = 32'h00008067;
mem['h0B47] = 32'h00000013;
mem['h0B48] = 32'h00812783;
mem['h0B49] = 32'h00178793;
mem['h0B4A] = 32'h00F12423;
mem['h0B4B] = 32'hF61FF06F;
mem['h0B4C] = 32'h96010113;
mem['h0B4D] = 32'h000065B7;
mem['h0B4E] = 32'h69412423;
mem['h0B4F] = 32'h02000613;
mem['h0B50] = 32'h9D858593;
mem['h0B51] = 32'h00050A13;
mem['h0B52] = 32'h03010513;
mem['h0B53] = 32'h68112E23;
mem['h0B54] = 32'h68812C23;
mem['h0B55] = 32'h68912A23;
mem['h0B56] = 32'h69212823;
mem['h0B57] = 32'h69312623;
mem['h0B58] = 32'h69612023;
mem['h0B59] = 32'h67712E23;
mem['h0B5A] = 32'h69512223;
mem['h0B5B] = 32'h895FF0EF;
mem['h0B5C] = 32'h000065B7;
mem['h0B5D] = 32'h00C00613;
mem['h0B5E] = 32'h77058593;
mem['h0B5F] = 32'h00410513;
mem['h0B60] = 32'h881FF0EF;
mem['h0B61] = 32'h00006B37;
mem['h0B62] = 32'h934B0513;
mem['h0B63] = 32'hF1CFD0EF;
mem['h0B64] = 32'h00006437;
mem['h0B65] = 32'h00050913;
mem['h0B66] = 32'h95440513;
mem['h0B67] = 32'hF0CFD0EF;
mem['h0B68] = 32'h00050493;
mem['h0B69] = 32'h00410613;
mem['h0B6A] = 32'h03010593;
mem['h0B6B] = 32'h17010513;
mem['h0B6C] = 32'hE09FF0EF;
mem['h0B6D] = 32'h95440593;
mem['h0B6E] = 32'h412009B3;
mem['h0B6F] = 32'h40900433;
mem['h0B70] = 32'h00048613;
mem['h0B71] = 32'h07010513;
mem['h0B72] = 32'h00100793;
mem['h0B73] = 32'h00410713;
mem['h0B74] = 32'h03010693;
mem['h0B75] = 32'h00F9F993;
mem['h0B76] = 32'h00F47413;
mem['h0B77] = 32'h849FF0EF;
mem['h0B78] = 32'h012989B3;
mem['h0B79] = 32'h00940433;
mem['h0B7A] = 32'h01340433;
mem['h0B7B] = 32'h40000613;
mem['h0B7C] = 32'h00000593;
mem['h0B7D] = 32'h27010513;
mem['h0B7E] = 32'h01040B93;
mem['h0B7F] = 32'hE20FF0EF;
mem['h0B80] = 32'h00090A63;
mem['h0B81] = 32'h00090613;
mem['h0B82] = 32'h934B0593;
mem['h0B83] = 32'h27010513;
mem['h0B84] = 32'hFF0FF0EF;
mem['h0B85] = 32'h27010793;
mem['h0B86] = 32'h00048613;
mem['h0B87] = 32'h07010593;
mem['h0B88] = 32'h01378533;
mem['h0B89] = 32'hFDCFF0EF;
mem['h0B8A] = 32'h27010793;
mem['h0B8B] = 32'h00878AB3;
mem['h0B8C] = 32'h00090593;
mem['h0B8D] = 32'h00000613;
mem['h0B8E] = 32'h000A8513;
mem['h0B8F] = 32'h851FD0EF;
mem['h0B90] = 32'h00048593;
mem['h0B91] = 32'h00000613;
mem['h0B92] = 32'h008A8513;
mem['h0B93] = 32'h841FD0EF;
mem['h0B94] = 32'h000B8693;
mem['h0B95] = 32'h27010613;
mem['h0B96] = 32'h17010593;
mem['h0B97] = 32'h01010513;
mem['h0B98] = 32'hB65FF0EF;
mem['h0B99] = 32'h00410613;
mem['h0B9A] = 32'h03010593;
mem['h0B9B] = 32'h05010513;
mem['h0B9C] = 32'hD49FF0EF;
mem['h0B9D] = 32'h40000613;
mem['h0B9E] = 32'h00000593;
mem['h0B9F] = 32'h27010513;
mem['h0BA0] = 32'hD9CFF0EF;
mem['h0BA1] = 32'h00090A63;
mem['h0BA2] = 32'h00090613;
mem['h0BA3] = 32'h934B0593;
mem['h0BA4] = 32'h27010513;
mem['h0BA5] = 32'hF6CFF0EF;
mem['h0BA6] = 32'h27010793;
mem['h0BA7] = 32'h00048613;
mem['h0BA8] = 32'h07010593;
mem['h0BA9] = 32'h01378533;
mem['h0BAA] = 32'hF58FF0EF;
mem['h0BAB] = 32'h27010793;
mem['h0BAC] = 32'h00878433;
mem['h0BAD] = 32'h00090593;
mem['h0BAE] = 32'h00000613;
mem['h0BAF] = 32'h00040513;
mem['h0BB0] = 32'hFCCFD0EF;
mem['h0BB1] = 32'h00048593;
mem['h0BB2] = 32'h00000613;
mem['h0BB3] = 32'h00840513;
mem['h0BB4] = 32'hFBCFD0EF;
mem['h0BB5] = 32'h000B8693;
mem['h0BB6] = 32'h27010613;
mem['h0BB7] = 32'h05010593;
mem['h0BB8] = 32'h02010513;
mem['h0BB9] = 32'hAE1FF0EF;
mem['h0BBA] = 32'h01012703;
mem['h0BBB] = 32'h02012783;
mem['h0BBC] = 32'h06F71E63;
mem['h0BBD] = 32'h01412703;
mem['h0BBE] = 32'h02412783;
mem['h0BBF] = 32'h06F71863;
mem['h0BC0] = 32'h01812703;
mem['h0BC1] = 32'h02812783;
mem['h0BC2] = 32'h06F71263;
mem['h0BC3] = 32'h01C12703;
mem['h0BC4] = 32'h02C12783;
mem['h0BC5] = 32'h04F71C63;
mem['h0BC6] = 32'h07010593;
mem['h0BC7] = 32'h00100793;
mem['h0BC8] = 32'h00410713;
mem['h0BC9] = 32'h03010693;
mem['h0BCA] = 32'h00048613;
mem['h0BCB] = 32'h17010513;
mem['h0BCC] = 32'hEF4FF0EF;
mem['h0BCD] = 32'h000065B7;
mem['h0BCE] = 32'h99058593;
mem['h0BCF] = 32'h69812403;
mem['h0BD0] = 32'h69C12083;
mem['h0BD1] = 32'h69412483;
mem['h0BD2] = 32'h69012903;
mem['h0BD3] = 32'h68C12983;
mem['h0BD4] = 32'h68412A83;
mem['h0BD5] = 32'h68012B03;
mem['h0BD6] = 32'h67C12B83;
mem['h0BD7] = 32'h000A0513;
mem['h0BD8] = 32'h68812A03;
mem['h0BD9] = 32'h6A010113;
mem['h0BDA] = 32'hA5CFD06F;
mem['h0BDB] = 32'h000065B7;
mem['h0BDC] = 32'h9B458593;
mem['h0BDD] = 32'hFC9FF06F;
mem['h0BDE] = 32'hE5010113;
mem['h0BDF] = 32'h03000513;
mem['h0BE0] = 32'h1A112623;
mem['h0BE1] = 32'h1A812423;
mem['h0BE2] = 32'h1A912223;
mem['h0BE3] = 32'h1B212023;
mem['h0BE4] = 32'h19312E23;
mem['h0BE5] = 32'h19412C23;
mem['h0BE6] = 32'h19512A23;
mem['h0BE7] = 32'h19612823;
mem['h0BE8] = 32'h19712623;
mem['h0BE9] = 32'h19812423;
mem['h0BEA] = 32'h19912223;
mem['h0BEB] = 32'h19A12023;
mem['h0BEC] = 32'h17B12E23;
mem['h0BED] = 32'h904FE0EF;
mem['h0BEE] = 32'h00050413;
mem['h0BEF] = 32'h00800513;
mem['h0BF0] = 32'h8F8FE0EF;
mem['h0BF1] = 32'h00050913;
mem['h0BF2] = 32'h01C00513;
mem['h0BF3] = 32'h8ECFE0EF;
mem['h0BF4] = 32'h00050493;
mem['h0BF5] = 32'h00400513;
mem['h0BF6] = 32'h8E0FE0EF;
mem['h0BF7] = 32'h200007B7;
mem['h0BF8] = 32'h00F52023;
mem['h0BF9] = 32'h00A4A023;
mem['h0BFA] = 32'h00400513;
mem['h0BFB] = 32'h8CCFE0EF;
mem['h0BFC] = 32'h200007B7;
mem['h0BFD] = 32'h00478793;
mem['h0BFE] = 32'h00F52023;
mem['h0BFF] = 32'h00A4A223;
mem['h0C00] = 32'h00400513;
mem['h0C01] = 32'h8B4FE0EF;
mem['h0C02] = 32'h200007B7;
mem['h0C03] = 32'h00878793;
mem['h0C04] = 32'h00F52023;
mem['h0C05] = 32'h00A4A423;
mem['h0C06] = 32'h00400513;
mem['h0C07] = 32'h89CFE0EF;
mem['h0C08] = 32'h200007B7;
mem['h0C09] = 32'h00C78793;
mem['h0C0A] = 32'h00F52023;
mem['h0C0B] = 32'h00A4A623;
mem['h0C0C] = 32'h00400513;
mem['h0C0D] = 32'h884FE0EF;
mem['h0C0E] = 32'h200007B7;
mem['h0C0F] = 32'h01078793;
mem['h0C10] = 32'h00F52023;
mem['h0C11] = 32'h00A4A823;
mem['h0C12] = 32'h00400513;
mem['h0C13] = 32'h86CFE0EF;
mem['h0C14] = 32'h200007B7;
mem['h0C15] = 32'h01478793;
mem['h0C16] = 32'h00F52023;
mem['h0C17] = 32'h00A4AA23;
mem['h0C18] = 32'h00400513;
mem['h0C19] = 32'h854FE0EF;
mem['h0C1A] = 32'h200007B7;
mem['h0C1B] = 32'h01878793;
mem['h0C1C] = 32'h00F52023;
mem['h0C1D] = 32'h00A4AC23;
mem['h0C1E] = 32'h00992023;
mem['h0C1F] = 32'h01C00513;
mem['h0C20] = 32'h838FE0EF;
mem['h0C21] = 32'h00050493;
mem['h0C22] = 32'h00400513;
mem['h0C23] = 32'h82CFE0EF;
mem['h0C24] = 32'h200007B7;
mem['h0C25] = 32'h01C78793;
mem['h0C26] = 32'h00F52023;
mem['h0C27] = 32'h00A4A023;
mem['h0C28] = 32'h00400513;
mem['h0C29] = 32'h814FE0EF;
mem['h0C2A] = 32'h200007B7;
mem['h0C2B] = 32'h02078793;
mem['h0C2C] = 32'h00F52023;
mem['h0C2D] = 32'h00A4A223;
mem['h0C2E] = 32'h00400513;
mem['h0C2F] = 32'hFFDFD0EF;
mem['h0C30] = 32'h200007B7;
mem['h0C31] = 32'h02478793;
mem['h0C32] = 32'h00F52023;
mem['h0C33] = 32'h00A4A423;
mem['h0C34] = 32'h00400513;
mem['h0C35] = 32'hFE5FD0EF;
mem['h0C36] = 32'h200007B7;
mem['h0C37] = 32'h02878793;
mem['h0C38] = 32'h00F52023;
mem['h0C39] = 32'h00A4A623;
mem['h0C3A] = 32'h00400513;
mem['h0C3B] = 32'hFCDFD0EF;
mem['h0C3C] = 32'h200007B7;
mem['h0C3D] = 32'h02C78793;
mem['h0C3E] = 32'h00F52023;
mem['h0C3F] = 32'h00A4A823;
mem['h0C40] = 32'h00400513;
mem['h0C41] = 32'hFB5FD0EF;
mem['h0C42] = 32'h200007B7;
mem['h0C43] = 32'h03078793;
mem['h0C44] = 32'h00F52023;
mem['h0C45] = 32'h00A4AA23;
mem['h0C46] = 32'h00400513;
mem['h0C47] = 32'hF9DFD0EF;
mem['h0C48] = 32'h200007B7;
mem['h0C49] = 32'h03478793;
mem['h0C4A] = 32'h00F52023;
mem['h0C4B] = 32'h00A4AC23;
mem['h0C4C] = 32'h00992223;
mem['h0C4D] = 32'h01242023;
mem['h0C4E] = 32'h01000513;
mem['h0C4F] = 32'hF7DFD0EF;
mem['h0C50] = 32'h00050493;
mem['h0C51] = 32'h00400513;
mem['h0C52] = 32'hF71FD0EF;
mem['h0C53] = 32'h200007B7;
mem['h0C54] = 32'h03878793;
mem['h0C55] = 32'h00F52023;
mem['h0C56] = 32'h00A4A023;
mem['h0C57] = 32'h00400513;
mem['h0C58] = 32'hF59FD0EF;
mem['h0C59] = 32'h200007B7;
mem['h0C5A] = 32'h03C78793;
mem['h0C5B] = 32'h00F52023;
mem['h0C5C] = 32'h00A4A223;
mem['h0C5D] = 32'h00400513;
mem['h0C5E] = 32'hF41FD0EF;
mem['h0C5F] = 32'h200007B7;
mem['h0C60] = 32'h04078793;
mem['h0C61] = 32'h00F52023;
mem['h0C62] = 32'h00A4A423;
mem['h0C63] = 32'h00400513;
mem['h0C64] = 32'hF29FD0EF;
mem['h0C65] = 32'h200007B7;
mem['h0C66] = 32'h04478793;
mem['h0C67] = 32'h00F52023;
mem['h0C68] = 32'h00A4A623;
mem['h0C69] = 32'h00942223;
mem['h0C6A] = 32'h00400513;
mem['h0C6B] = 32'hF0DFD0EF;
mem['h0C6C] = 32'h200007B7;
mem['h0C6D] = 32'h04878793;
mem['h0C6E] = 32'h00F52023;
mem['h0C6F] = 32'h200004B7;
mem['h0C70] = 32'h200009B7;
mem['h0C71] = 32'h00A42423;
mem['h0C72] = 32'h00C40A13;
mem['h0C73] = 32'h04C48493;
mem['h0C74] = 32'h07C98993;
mem['h0C75] = 32'h00C00513;
mem['h0C76] = 32'hEE1FD0EF;
mem['h0C77] = 32'h00050913;
mem['h0C78] = 32'h00400513;
mem['h0C79] = 32'hED5FD0EF;
mem['h0C7A] = 32'h00952023;
mem['h0C7B] = 32'h00A92023;
mem['h0C7C] = 32'h00400513;
mem['h0C7D] = 32'hEC5FD0EF;
mem['h0C7E] = 32'h00448793;
mem['h0C7F] = 32'h00F52023;
mem['h0C80] = 32'h00A92223;
mem['h0C81] = 32'h00400513;
mem['h0C82] = 32'hEB1FD0EF;
mem['h0C83] = 32'h00848793;
mem['h0C84] = 32'h00F52023;
mem['h0C85] = 32'h00A92423;
mem['h0C86] = 32'h012A2023;
mem['h0C87] = 32'h00C48493;
mem['h0C88] = 32'h004A0A13;
mem['h0C89] = 32'hFB3498E3;
mem['h0C8A] = 32'h00400513;
mem['h0C8B] = 32'hE8DFD0EF;
mem['h0C8C] = 32'h00952023;
mem['h0C8D] = 32'h00A42E23;
mem['h0C8E] = 32'h00400513;
mem['h0C8F] = 32'hE7DFD0EF;
mem['h0C90] = 32'h200007B7;
mem['h0C91] = 32'h08078793;
mem['h0C92] = 32'h00F52023;
mem['h0C93] = 32'h02A42023;
mem['h0C94] = 32'h00400513;
mem['h0C95] = 32'hE65FD0EF;
mem['h0C96] = 32'h00050493;
mem['h0C97] = 32'h00400513;
mem['h0C98] = 32'hE59FD0EF;
mem['h0C99] = 32'h200007B7;
mem['h0C9A] = 32'h08478793;
mem['h0C9B] = 32'h00F52023;
mem['h0C9C] = 32'h00A4A023;
mem['h0C9D] = 32'h02942223;
mem['h0C9E] = 32'h10000513;
mem['h0C9F] = 32'hE3DFD0EF;
mem['h0CA0] = 32'h200004B7;
mem['h0CA1] = 32'h20001A37;
mem['h0CA2] = 32'h00050913;
mem['h0CA3] = 32'h00050A93;
mem['h0CA4] = 32'h40048493;
mem['h0CA5] = 32'h800A0A13;
mem['h0CA6] = 32'h01000513;
mem['h0CA7] = 32'hE1DFD0EF;
mem['h0CA8] = 32'h00050993;
mem['h0CA9] = 32'h00400513;
mem['h0CAA] = 32'hE11FD0EF;
mem['h0CAB] = 32'h00952023;
mem['h0CAC] = 32'h00A9A023;
mem['h0CAD] = 32'h00400513;
mem['h0CAE] = 32'hE01FD0EF;
mem['h0CAF] = 32'h00448793;
mem['h0CB0] = 32'h00F52023;
mem['h0CB1] = 32'h00A9A223;
mem['h0CB2] = 32'h00400513;
mem['h0CB3] = 32'hDEDFD0EF;
mem['h0CB4] = 32'h00848793;
mem['h0CB5] = 32'h00F52023;
mem['h0CB6] = 32'h00A9A423;
mem['h0CB7] = 32'h00400513;
mem['h0CB8] = 32'hDD9FD0EF;
mem['h0CB9] = 32'h00C48793;
mem['h0CBA] = 32'h00F52023;
mem['h0CBB] = 32'h00A9A623;
mem['h0CBC] = 32'h013AA023;
mem['h0CBD] = 32'h01048493;
mem['h0CBE] = 32'h004A8A93;
mem['h0CBF] = 32'hF9449EE3;
mem['h0CC0] = 32'h03242423;
mem['h0CC1] = 32'h10000513;
mem['h0CC2] = 32'hDB1FD0EF;
mem['h0CC3] = 32'h20004A37;
mem['h0CC4] = 32'h00050993;
mem['h0CC5] = 32'h00050A93;
mem['h0CC6] = 32'h200024B7;
mem['h0CC7] = 32'hE00A0A13;
mem['h0CC8] = 32'h07800513;
mem['h0CC9] = 32'hD95FD0EF;
mem['h0CCA] = 32'h00050913;
mem['h0CCB] = 32'h00400513;
mem['h0CCC] = 32'hD89FD0EF;
mem['h0CCD] = 32'h00952023;
mem['h0CCE] = 32'h00A92023;
mem['h0CCF] = 32'h00400513;
mem['h0CD0] = 32'hD79FD0EF;
mem['h0CD1] = 32'h00448793;
mem['h0CD2] = 32'h00F52023;
mem['h0CD3] = 32'h00A92223;
mem['h0CD4] = 32'h00400513;
mem['h0CD5] = 32'hD65FD0EF;
mem['h0CD6] = 32'h00848793;
mem['h0CD7] = 32'h00F52023;
mem['h0CD8] = 32'h00A92423;
mem['h0CD9] = 32'h00400513;
mem['h0CDA] = 32'hD51FD0EF;
mem['h0CDB] = 32'h00C48793;
mem['h0CDC] = 32'h00F52023;
mem['h0CDD] = 32'h00A92623;
mem['h0CDE] = 32'h00400513;
mem['h0CDF] = 32'hD3DFD0EF;
mem['h0CE0] = 32'h01048793;
mem['h0CE1] = 32'h00F52023;
mem['h0CE2] = 32'h00A92823;
mem['h0CE3] = 32'h00400513;
mem['h0CE4] = 32'hD29FD0EF;
mem['h0CE5] = 32'h01448793;
mem['h0CE6] = 32'h00F52023;
mem['h0CE7] = 32'h00A92A23;
mem['h0CE8] = 32'h00400513;
mem['h0CE9] = 32'hD15FD0EF;
mem['h0CEA] = 32'h01848793;
mem['h0CEB] = 32'h00F52023;
mem['h0CEC] = 32'h00A92C23;
mem['h0CED] = 32'h00400513;
mem['h0CEE] = 32'hD01FD0EF;
mem['h0CEF] = 32'h01C48793;
mem['h0CF0] = 32'h00F52023;
mem['h0CF1] = 32'h00A92E23;
mem['h0CF2] = 32'h00400513;
mem['h0CF3] = 32'hCEDFD0EF;
mem['h0CF4] = 32'h02048793;
mem['h0CF5] = 32'h00F52023;
mem['h0CF6] = 32'h02A92023;
mem['h0CF7] = 32'h00400513;
mem['h0CF8] = 32'hCD9FD0EF;
mem['h0CF9] = 32'h02448793;
mem['h0CFA] = 32'h00F52023;
mem['h0CFB] = 32'h02A92223;
mem['h0CFC] = 32'h00400513;
mem['h0CFD] = 32'hCC5FD0EF;
mem['h0CFE] = 32'h02848793;
mem['h0CFF] = 32'h00F52023;
mem['h0D00] = 32'h02A92423;
mem['h0D01] = 32'h00400513;
mem['h0D02] = 32'hCB1FD0EF;
mem['h0D03] = 32'h02C48793;
mem['h0D04] = 32'h00F52023;
mem['h0D05] = 32'h02A92623;
mem['h0D06] = 32'h00400513;
mem['h0D07] = 32'hC9DFD0EF;
mem['h0D08] = 32'h03048793;
mem['h0D09] = 32'h00F52023;
mem['h0D0A] = 32'h02A92823;
mem['h0D0B] = 32'h00400513;
mem['h0D0C] = 32'hC89FD0EF;
mem['h0D0D] = 32'h03448793;
mem['h0D0E] = 32'h00F52023;
mem['h0D0F] = 32'h02A92A23;
mem['h0D10] = 32'h00400513;
mem['h0D11] = 32'hC75FD0EF;
mem['h0D12] = 32'h03848793;
mem['h0D13] = 32'h00F52023;
mem['h0D14] = 32'h02A92C23;
mem['h0D15] = 32'h00400513;
mem['h0D16] = 32'hC61FD0EF;
mem['h0D17] = 32'h03C48793;
mem['h0D18] = 32'h00F52023;
mem['h0D19] = 32'h02A92E23;
mem['h0D1A] = 32'h00400513;
mem['h0D1B] = 32'hC4DFD0EF;
mem['h0D1C] = 32'h04048793;
mem['h0D1D] = 32'h00F52023;
mem['h0D1E] = 32'h04A92023;
mem['h0D1F] = 32'h00400513;
mem['h0D20] = 32'hC39FD0EF;
mem['h0D21] = 32'h04448793;
mem['h0D22] = 32'h00F52023;
mem['h0D23] = 32'h04A92223;
mem['h0D24] = 32'h00400513;
mem['h0D25] = 32'hC25FD0EF;
mem['h0D26] = 32'h04848793;
mem['h0D27] = 32'h00F52023;
mem['h0D28] = 32'h04A92423;
mem['h0D29] = 32'h00400513;
mem['h0D2A] = 32'hC11FD0EF;
mem['h0D2B] = 32'h04C48793;
mem['h0D2C] = 32'h00F52023;
mem['h0D2D] = 32'h04A92623;
mem['h0D2E] = 32'h00400513;
mem['h0D2F] = 32'hBFDFD0EF;
mem['h0D30] = 32'h05048793;
mem['h0D31] = 32'h00F52023;
mem['h0D32] = 32'h04A92823;
mem['h0D33] = 32'h00400513;
mem['h0D34] = 32'hBE9FD0EF;
mem['h0D35] = 32'h05448793;
mem['h0D36] = 32'h00F52023;
mem['h0D37] = 32'h04A92A23;
mem['h0D38] = 32'h00400513;
mem['h0D39] = 32'hBD5FD0EF;
mem['h0D3A] = 32'h05848793;
mem['h0D3B] = 32'h00F52023;
mem['h0D3C] = 32'h04A92C23;
mem['h0D3D] = 32'h00400513;
mem['h0D3E] = 32'hBC1FD0EF;
mem['h0D3F] = 32'h05C48793;
mem['h0D40] = 32'h00F52023;
mem['h0D41] = 32'h04A92E23;
mem['h0D42] = 32'h00400513;
mem['h0D43] = 32'hBADFD0EF;
mem['h0D44] = 32'h06048793;
mem['h0D45] = 32'h00F52023;
mem['h0D46] = 32'h06A92023;
mem['h0D47] = 32'h00400513;
mem['h0D48] = 32'hB99FD0EF;
mem['h0D49] = 32'h06448793;
mem['h0D4A] = 32'h00F52023;
mem['h0D4B] = 32'h06A92223;
mem['h0D4C] = 32'h00400513;
mem['h0D4D] = 32'hB85FD0EF;
mem['h0D4E] = 32'h06848793;
mem['h0D4F] = 32'h00F52023;
mem['h0D50] = 32'h06A92423;
mem['h0D51] = 32'h00400513;
mem['h0D52] = 32'hB71FD0EF;
mem['h0D53] = 32'h06C48793;
mem['h0D54] = 32'h00F52023;
mem['h0D55] = 32'h06A92623;
mem['h0D56] = 32'h00400513;
mem['h0D57] = 32'hB5DFD0EF;
mem['h0D58] = 32'h07048793;
mem['h0D59] = 32'h00F52023;
mem['h0D5A] = 32'h06A92823;
mem['h0D5B] = 32'h00400513;
mem['h0D5C] = 32'hB49FD0EF;
mem['h0D5D] = 32'h07448793;
mem['h0D5E] = 32'h00F52023;
mem['h0D5F] = 32'h06A92A23;
mem['h0D60] = 32'h012AA023;
mem['h0D61] = 32'h07848493;
mem['h0D62] = 32'h004A8A93;
mem['h0D63] = 32'hD9449AE3;
mem['h0D64] = 32'h01C42783;
mem['h0D65] = 32'h03342623;
mem['h0D66] = 32'h0007A783;
mem['h0D67] = 32'h0027D703;
mem['h0D68] = 32'h0000D7B7;
mem['h0D69] = 32'hCBA78793;
mem['h0D6A] = 32'h00F71E63;
mem['h0D6B] = 32'h01C42783;
mem['h0D6C] = 32'h0007A783;
mem['h0D6D] = 32'h0007D703;
mem['h0D6E] = 32'h0000D7B7;
mem['h0D6F] = 32'hACA78793;
mem['h0D70] = 32'h00F70C63;
mem['h0D71] = 32'h000065B7;
mem['h0D72] = 32'h9FC58593;
mem['h0D73] = 32'h00040513;
mem['h0D74] = 32'hBF5FC0EF;
mem['h0D75] = 32'h00100073;
mem['h0D76] = 32'h000065B7;
mem['h0D77] = 32'hA2458593;
mem['h0D78] = 32'h00040513;
mem['h0D79] = 32'hBE1FC0EF;
mem['h0D7A] = 32'h000065B7;
mem['h0D7B] = 32'hA5458593;
mem['h0D7C] = 32'h00040513;
mem['h0D7D] = 32'hBD1FC0EF;
mem['h0D7E] = 32'h02042783;
mem['h0D7F] = 32'h00040513;
mem['h0D80] = 32'h100009B7;
mem['h0D81] = 32'h0007A783;
mem['h0D82] = 32'h00098493;
mem['h0D83] = 32'h0037C583;
mem['h0D84] = 32'hAF9FC0EF;
mem['h0D85] = 32'h02E00593;
mem['h0D86] = 32'h00040513;
mem['h0D87] = 32'hA59FC0EF;
mem['h0D88] = 32'h02042783;
mem['h0D89] = 32'h00040513;
mem['h0D8A] = 32'h0007A783;
mem['h0D8B] = 32'h0027C583;
mem['h0D8C] = 32'hAD9FC0EF;
mem['h0D8D] = 32'h02E00593;
mem['h0D8E] = 32'h00040513;
mem['h0D8F] = 32'hA39FC0EF;
mem['h0D90] = 32'h02042783;
mem['h0D91] = 32'h00040513;
mem['h0D92] = 32'h0007A783;
mem['h0D93] = 32'h0007D583;
mem['h0D94] = 32'hAB9FC0EF;
mem['h0D95] = 32'h000065B7;
mem['h0D96] = 32'hA7058593;
mem['h0D97] = 32'h00040513;
mem['h0D98] = 32'hB65FC0EF;
mem['h0D99] = 32'h000065B7;
mem['h0D9A] = 32'hAA058593;
mem['h0D9B] = 32'h00040513;
mem['h0D9C] = 32'hB55FC0EF;
mem['h0D9D] = 32'h000065B7;
mem['h0D9E] = 32'hAD058593;
mem['h0D9F] = 32'h00040513;
mem['h0DA0] = 32'hB45FC0EF;
mem['h0DA1] = 32'h00098713;
mem['h0DA2] = 32'h00174683;
mem['h0DA3] = 32'h00074783;
mem['h0DA4] = 32'h00D7E7B3;
mem['h0DA5] = 32'h00274683;
mem['h0DA6] = 32'h00374703;
mem['h0DA7] = 32'h00D7E7B3;
mem['h0DA8] = 32'h00E7E7B3;
mem['h0DA9] = 32'h04079263;
mem['h0DAA] = 32'h6201B7B7;
mem['h0DAB] = 32'h8C078793;
mem['h0DAC] = 32'h00F4A023;
mem['h0DAD] = 32'h010007B7;
mem['h0DAE] = 32'hFFF78793;
mem['h0DAF] = 32'h00F4A223;
mem['h0DB0] = 32'hCACAC7B7;
mem['h0DB1] = 32'hACC78793;
mem['h0DB2] = 32'h00F4A423;
mem['h0DB3] = 32'hA8C007B7;
mem['h0DB4] = 32'h10078793;
mem['h0DB5] = 32'h00F4A623;
mem['h0DB6] = 32'hE0100793;
mem['h0DB7] = 32'h00F49823;
mem['h0DB8] = 32'h00100793;
mem['h0DB9] = 32'h00F48923;
mem['h0DBA] = 32'h00040513;
mem['h0DBB] = 32'h904FE0EF;
mem['h0DBC] = 32'h000065B7;
mem['h0DBD] = 32'hAE058593;
mem['h0DBE] = 32'h00040513;
mem['h0DBF] = 32'hAC9FC0EF;
mem['h0DC0] = 32'h00006BB7;
mem['h0DC1] = 32'hB08B8593;
mem['h0DC2] = 32'h00040513;
mem['h0DC3] = 32'hAB9FC0EF;
mem['h0DC4] = 32'h81418793;
mem['h0DC5] = 32'h00F12023;
mem['h0DC6] = 32'h00006AB7;
mem['h0DC7] = 32'h61C48793;
mem['h0DC8] = 32'h00000913;
mem['h0DC9] = 32'h00F12223;
mem['h0DCA] = 32'h630A8A93;
mem['h0DCB] = 32'h5F000C13;
mem['h0DCC] = 32'h60000C93;
mem['h0DCD] = 32'h00800D13;
mem['h0DCE] = 32'h00100B13;
mem['h0DCF] = 32'h00200D93;
mem['h0DD0] = 32'h00048A23;
mem['h0DD1] = 32'h00049B23;
mem['h0DD2] = 32'h00042783;
mem['h0DD3] = 32'h0047A783;
mem['h0DD4] = 32'h0187A783;
mem['h0DD5] = 32'h0007A783;
mem['h0DD6] = 32'h0007A783;
mem['h0DD7] = 32'h0017F793;
mem['h0DD8] = 32'h0E078E63;
mem['h0DD9] = 32'h00042783;
mem['h0DDA] = 32'h01448713;
mem['h0DDB] = 32'h0047A783;
mem['h0DDC] = 32'h0107A783;
mem['h0DDD] = 32'h0007A783;
mem['h0DDE] = 32'h0007A783;
mem['h0DDF] = 32'h0037D793;
mem['h0DE0] = 32'h0077F793;
mem['h0DE1] = 32'h00F48AA3;
mem['h0DE2] = 32'h00000793;
mem['h0DE3] = 32'h06FC6263;
mem['h0DE4] = 32'h00042683;
mem['h0DE5] = 32'h0046A683;
mem['h0DE6] = 32'h0006A683;
mem['h0DE7] = 32'h0006A683;
mem['h0DE8] = 32'h0006A683;
mem['h0DE9] = 32'h00D72423;
mem['h0DEA] = 32'h00042683;
mem['h0DEB] = 32'h0046A683;
mem['h0DEC] = 32'h0046A683;
mem['h0DED] = 32'h0006A683;
mem['h0DEE] = 32'h0006A683;
mem['h0DEF] = 32'h00D72623;
mem['h0DF0] = 32'h00042683;
mem['h0DF1] = 32'h0046A683;
mem['h0DF2] = 32'h0086A683;
mem['h0DF3] = 32'h0006A683;
mem['h0DF4] = 32'h0006A683;
mem['h0DF5] = 32'h00D72823;
mem['h0DF6] = 32'h00042683;
mem['h0DF7] = 32'h0046A683;
mem['h0DF8] = 32'h00C6A683;
mem['h0DF9] = 32'h0006A683;
mem['h0DFA] = 32'h0006A683;
mem['h0DFB] = 32'h00D72A23;
mem['h0DFC] = 32'h00042683;
mem['h0DFD] = 32'h01070713;
mem['h0DFE] = 32'h0046A683;
mem['h0DFF] = 32'h0106A683;
mem['h0E00] = 32'h0006A683;
mem['h0E01] = 32'h0006A683;
mem['h0E02] = 32'h01069613;
mem['h0E03] = 32'h06065A63;
mem['h0E04] = 32'h00042703;
mem['h0E05] = 32'h00472703;
mem['h0E06] = 32'h01072703;
mem['h0E07] = 32'h00072703;
mem['h0E08] = 32'h00275703;
mem['h0E09] = 32'h00177693;
mem['h0E0A] = 32'h04069663;
mem['h0E0B] = 32'h00FCF463;
mem['h0E0C] = 32'h60000793;
mem['h0E0D] = 32'h00F4AC23;
mem['h0E0E] = 32'h00042783;
mem['h0E0F] = 32'h0047A783;
mem['h0E10] = 32'h0147A783;
mem['h0E11] = 32'h0007A703;
mem['h0E12] = 32'h00072783;
mem['h0E13] = 32'h0017E793;
mem['h0E14] = 32'h00F72023;
mem['h0E15] = 32'h0184A783;
mem['h0E16] = 32'h04079663;
mem['h0E17] = 32'h00842783;
mem['h0E18] = 32'h0007A703;
mem['h0E19] = 32'h00072783;
mem['h0E1A] = 32'hDFF7F793;
mem['h0E1B] = 32'h00F72023;
mem['h0E1C] = 32'h3580006F;
mem['h0E1D] = 32'h00178793;
mem['h0E1E] = 32'h00175713;
mem['h0E1F] = 32'hFA9FF06F;
mem['h0E20] = 32'h00042683;
mem['h0E21] = 32'h01078793;
mem['h0E22] = 32'h0046A683;
mem['h0E23] = 32'h0146A683;
mem['h0E24] = 32'h0006A603;
mem['h0E25] = 32'h00062683;
mem['h0E26] = 32'h0016E693;
mem['h0E27] = 32'h00D62023;
mem['h0E28] = 32'hEEDFF06F;
mem['h0E29] = 32'h00842783;
mem['h0E2A] = 32'h0007A703;
mem['h0E2B] = 32'h00072783;
mem['h0E2C] = 32'h2007E793;
mem['h0E2D] = 32'h00F72023;
mem['h0E2E] = 32'h0284C783;
mem['h0E2F] = 32'h35A79663;
mem['h0E30] = 32'h0294C783;
mem['h0E31] = 32'h00600713;
mem['h0E32] = 32'h18E78663;
mem['h0E33] = 32'h32079E63;
mem['h0E34] = 32'h02A4C783;
mem['h0E35] = 32'h04000713;
mem['h0E36] = 32'h0F07F793;
mem['h0E37] = 32'h32E79663;
mem['h0E38] = 32'h0334C783;
mem['h0E39] = 32'h00100713;
mem['h0E3A] = 32'h00E78E63;
mem['h0E3B] = 32'h01100713;
mem['h0E3C] = 32'h30E79C63;
mem['h0E3D] = 32'h2A090A63;
mem['h0E3E] = 32'h000065B7;
mem['h0E3F] = 32'hB8458593;
mem['h0E40] = 32'h3140006F;
mem['h0E41] = 32'h02090863;
mem['h0E42] = 32'h000065B7;
mem['h0E43] = 32'hB5C58593;
mem['h0E44] = 32'h00040513;
mem['h0E45] = 32'h8B1FC0EF;
mem['h0E46] = 32'h0184A583;
mem['h0E47] = 32'h00040513;
mem['h0E48] = 32'hFE8FC0EF;
mem['h0E49] = 32'h000065B7;
mem['h0E4A] = 32'hBF058593;
mem['h0E4B] = 32'h00040513;
mem['h0E4C] = 32'h895FC0EF;
mem['h0E4D] = 32'h00400613;
mem['h0E4E] = 32'h00098593;
mem['h0E4F] = 32'h03A48513;
mem['h0E50] = 32'hB35FC0EF;
mem['h0E51] = 32'h0154C783;
mem['h0E52] = 32'h26051063;
mem['h0E53] = 32'h03E4C683;
mem['h0E54] = 32'h00800713;
mem['h0E55] = 32'h24E69A63;
mem['h0E56] = 32'h03F4C703;
mem['h0E57] = 32'h24071663;
mem['h0E58] = 32'h0184AA03;
mem['h0E59] = 32'h60F48E23;
mem['h0E5A] = 32'h00600613;
mem['h0E5B] = 32'h00100793;
mem['h0E5C] = 32'h02248593;
mem['h0E5D] = 32'h62448513;
mem['h0E5E] = 32'h60F48FA3;
mem['h0E5F] = 32'h6344A023;
mem['h0E60] = 32'hC81FE0EF;
mem['h0E61] = 32'h00600613;
mem['h0E62] = 32'h00848593;
mem['h0E63] = 32'h62A48513;
mem['h0E64] = 32'hC71FE0EF;
mem['h0E65] = 32'h00450737;
mem['h0E66] = 32'h00870713;
mem['h0E67] = 32'h62E4A823;
mem['h0E68] = 32'h02C4D703;
mem['h0E69] = 32'h00400613;
mem['h0E6A] = 32'h00098593;
mem['h0E6B] = 32'h62E49A23;
mem['h0E6C] = 32'h63E48513;
mem['h0E6D] = 32'h01FF0737;
mem['h0E6E] = 32'h62E4AC23;
mem['h0E6F] = 32'h62049B23;
mem['h0E70] = 32'h62049E23;
mem['h0E71] = 32'hC3DFE0EF;
mem['h0E72] = 32'h00400613;
mem['h0E73] = 32'h03648593;
mem['h0E74] = 32'h64248513;
mem['h0E75] = 32'hC2DFE0EF;
mem['h0E76] = 32'h01400593;
mem['h0E77] = 32'h63248513;
mem['h0E78] = 32'hA09FC0EF;
mem['h0E79] = 32'h00851713;
mem['h0E7A] = 32'h00855513;
mem['h0E7B] = 32'h00A76733;
mem['h0E7C] = 32'h62E49E23;
mem['h0E7D] = 32'h0424D703;
mem['h0E7E] = 32'hFD6A0613;
mem['h0E7F] = 32'h04648593;
mem['h0E80] = 32'h64E49523;
mem['h0E81] = 32'h0444D703;
mem['h0E82] = 32'h64E48513;
mem['h0E83] = 32'h64049323;
mem['h0E84] = 32'h64E49623;
mem['h0E85] = 32'h64049423;
mem['h0E86] = 32'hBE9FE0EF;
mem['h0E87] = 32'hFDEA0593;
mem['h0E88] = 32'h64648513;
mem['h0E89] = 32'h9C5FC0EF;
mem['h0E8A] = 32'h00851793;
mem['h0E8B] = 32'h00855513;
mem['h0E8C] = 32'h00A7E7B3;
mem['h0E8D] = 32'h64F49423;
mem['h0E8E] = 32'hE1C18593;
mem['h0E8F] = 32'h00040513;
mem['h0E90] = 32'hDECFE0EF;
mem['h0E91] = 32'h16090263;
mem['h0E92] = 32'h000065B7;
mem['h0E93] = 32'hB7058593;
mem['h0E94] = 32'h1340006F;
mem['h0E95] = 32'h02090863;
mem['h0E96] = 32'h000065B7;
mem['h0E97] = 32'hB3458593;
mem['h0E98] = 32'h00040513;
mem['h0E99] = 32'hF60FC0EF;
mem['h0E9A] = 32'h0184A583;
mem['h0E9B] = 32'h00040513;
mem['h0E9C] = 32'hE98FC0EF;
mem['h0E9D] = 32'h000065B7;
mem['h0E9E] = 32'hBF058593;
mem['h0E9F] = 32'h00040513;
mem['h0EA0] = 32'hF44FC0EF;
mem['h0EA1] = 32'h0154C703;
mem['h0EA2] = 32'h02B4CA03;
mem['h0EA3] = 32'h00100693;
mem['h0EA4] = 32'h00E12423;
mem['h0EA5] = 32'h02A4C783;
mem['h0EA6] = 32'h10DA1863;
mem['h0EA7] = 32'h02C4C603;
mem['h0EA8] = 32'h00800693;
mem['h0EA9] = 32'h10D61263;
mem['h0EAA] = 32'h02D4C683;
mem['h0EAB] = 32'h00D7E7B3;
mem['h0EAC] = 32'h0E079C63;
mem['h0EAD] = 32'h00400613;
mem['h0EAE] = 32'h00098593;
mem['h0EAF] = 32'h04248513;
mem['h0EB0] = 32'h9B5FC0EF;
mem['h0EB1] = 32'h0E051263;
mem['h0EB2] = 32'h0304C783;
mem['h0EB3] = 32'h0C079E63;
mem['h0EB4] = 32'h0314C783;
mem['h0EB5] = 32'h00812703;
mem['h0EB6] = 32'h0D479863;
mem['h0EB7] = 32'h60F48FA3;
mem['h0EB8] = 32'h00600613;
mem['h0EB9] = 32'h02A00793;
mem['h0EBA] = 32'h83218593;
mem['h0EBB] = 32'h62448513;
mem['h0EBC] = 32'h60E48E23;
mem['h0EBD] = 32'h62F4A023;
mem['h0EBE] = 32'hB09FE0EF;
mem['h0EBF] = 32'h00848593;
mem['h0EC0] = 32'h00600613;
mem['h0EC1] = 32'h62A48513;
mem['h0EC2] = 32'hAF9FE0EF;
mem['h0EC3] = 32'h010007B7;
mem['h0EC4] = 32'h60878793;
mem['h0EC5] = 32'h62F4A823;
mem['h0EC6] = 32'h040607B7;
mem['h0EC7] = 32'h00878793;
mem['h0EC8] = 32'h62F4AA23;
mem['h0EC9] = 32'h20000793;
mem['h0ECA] = 32'h62F49C23;
mem['h0ECB] = 32'h80818593;
mem['h0ECC] = 32'h00600613;
mem['h0ECD] = 32'h63A48513;
mem['h0ECE] = 32'hAC9FE0EF;
mem['h0ECF] = 32'h00400613;
mem['h0ED0] = 32'h00098593;
mem['h0ED1] = 32'h64048513;
mem['h0ED2] = 32'hAB9FE0EF;
mem['h0ED3] = 32'h00600613;
mem['h0ED4] = 32'h83218593;
mem['h0ED5] = 32'h64448513;
mem['h0ED6] = 32'hAA9FE0EF;
mem['h0ED7] = 32'h03848593;
mem['h0ED8] = 32'h00400613;
mem['h0ED9] = 32'h64A48513;
mem['h0EDA] = 32'hA99FE0EF;
mem['h0EDB] = 32'h00412583;
mem['h0EDC] = 32'h00040513;
mem['h0EDD] = 32'hCB8FE0EF;
mem['h0EDE] = 32'h02090863;
mem['h0EDF] = 32'h000065B7;
mem['h0EE0] = 32'hB4858593;
mem['h0EE1] = 32'h00040513;
mem['h0EE2] = 32'hE3CFC0EF;
mem['h0EE3] = 32'h6204A583;
mem['h0EE4] = 32'h00040513;
mem['h0EE5] = 32'hD74FC0EF;
mem['h0EE6] = 32'h000065B7;
mem['h0EE7] = 32'hBF058593;
mem['h0EE8] = 32'h00040513;
mem['h0EE9] = 32'hE20FC0EF;
mem['h0EEA] = 32'h0154C783;
mem['h0EEB] = 32'h07679C63;
mem['h0EEC] = 32'h00200793;
mem['h0EED] = 32'h00F48A23;
mem['h0EEE] = 32'h00012583;
mem['h0EEF] = 32'h00040513;
mem['h0EF0] = 32'h01648BA3;
mem['h0EF1] = 32'hC68FE0EF;
mem['h0EF2] = 32'h06810593;
mem['h0EF3] = 32'h00040513;
mem['h0EF4] = 32'hEB0FC0EF;
mem['h0EF5] = 32'h00050A13;
mem['h0EF6] = 32'hB60504E3;
mem['h0EF7] = 32'h000065B7;
mem['h0EF8] = 32'hB9858593;
mem['h0EF9] = 32'h06810513;
mem['h0EFA] = 32'h8E1FC0EF;
mem['h0EFB] = 32'h04051263;
mem['h0EFC] = 32'h00040513;
mem['h0EFD] = 32'h93CFF0EF;
mem['h0EFE] = 32'hB08B8593;
mem['h0EFF] = 32'h00040513;
mem['h0F00] = 32'hDC4FC0EF;
mem['h0F01] = 32'hB29FF06F;
mem['h0F02] = 32'hFA0900E3;
mem['h0F03] = 32'h000067B7;
mem['h0F04] = 32'hB1C78593;
mem['h0F05] = 32'h00040513;
mem['h0F06] = 32'hDACFC0EF;
mem['h0F07] = 32'h0184A583;
mem['h0F08] = 32'hF71FF06F;
mem['h0F09] = 32'hFBB792E3;
mem['h0F0A] = 32'h01648A23;
mem['h0F0B] = 32'hF8DFF06F;
mem['h0F0C] = 32'h000065B7;
mem['h0F0D] = 32'hBB058593;
mem['h0F0E] = 32'h06810513;
mem['h0F0F] = 32'h88DFC0EF;
mem['h0F10] = 32'h00050B13;
mem['h0F11] = 32'h0C051863;
mem['h0F12] = 32'h04800613;
mem['h0F13] = 32'h14CA8593;
mem['h0F14] = 32'h12810513;
mem['h0F15] = 32'h9ADFE0EF;
mem['h0F16] = 32'h00006A37;
mem['h0F17] = 32'h9D4A0513;
mem['h0F18] = 32'h849FC0EF;
mem['h0F19] = 32'h00050613;
mem['h0F1A] = 32'h9D4A0593;
mem['h0F1B] = 32'h10810513;
mem['h0F1C] = 32'hDD4FE0EF;
mem['h0F1D] = 32'h12810A13;
mem['h0F1E] = 32'h000A0713;
mem['h0F1F] = 32'h00000793;
mem['h0F20] = 32'h02000613;
mem['h0F21] = 32'h10810693;
mem['h0F22] = 32'h00F686B3;
mem['h0F23] = 32'h00474583;
mem['h0F24] = 32'h0006C683;
mem['h0F25] = 32'h06D59263;
mem['h0F26] = 32'h00178793;
mem['h0F27] = 32'h00170713;
mem['h0F28] = 32'hFEC792E3;
mem['h0F29] = 32'h00100C13;
mem['h0F2A] = 32'h00006CB7;
mem['h0F2B] = 32'hBC0C8513;
mem['h0F2C] = 32'hFF8FC0EF;
mem['h0F2D] = 32'h00050613;
mem['h0F2E] = 32'hBC0C8593;
mem['h0F2F] = 32'h10810513;
mem['h0F30] = 32'hD84FE0EF;
mem['h0F31] = 32'h02000793;
mem['h0F32] = 32'h10810713;
mem['h0F33] = 32'h01670733;
mem['h0F34] = 32'h00074683;
mem['h0F35] = 32'h028A4703;
mem['h0F36] = 32'h00E69A63;
mem['h0F37] = 32'h001B0B13;
mem['h0F38] = 32'h001A0A13;
mem['h0F39] = 32'hFEFB12E3;
mem['h0F3A] = 32'h000C1C63;
mem['h0F3B] = 32'h000065B7;
mem['h0F3C] = 32'hBDC58593;
mem['h0F3D] = 32'h0140006F;
mem['h0F3E] = 32'h00000C13;
mem['h0F3F] = 32'hFADFF06F;
mem['h0F40] = 32'h000065B7;
mem['h0F41] = 32'hBC458593;
mem['h0F42] = 32'h00040513;
mem['h0F43] = 32'hCB8FC0EF;
mem['h0F44] = 32'hEE9FF06F;
mem['h0F45] = 32'h000065B7;
mem['h0F46] = 32'hBF458593;
mem['h0F47] = 32'h06810513;
mem['h0F48] = 32'hFA8FC0EF;
mem['h0F49] = 32'h08051263;
mem['h0F4A] = 32'h08810513;
mem['h0F4B] = 32'hEF1FE0EF;
mem['h0F4C] = 32'h0A810513;
mem['h0F4D] = 32'hEE9FE0EF;
mem['h0F4E] = 32'h00006A37;
mem['h0F4F] = 32'h7C4A0613;
mem['h0F50] = 32'h08810593;
mem['h0F51] = 32'h0C810513;
mem['h0F52] = 32'hC99FD0EF;
mem['h0F53] = 32'h7C4A0613;
mem['h0F54] = 32'h0A810593;
mem['h0F55] = 32'h0E810513;
mem['h0F56] = 32'hC89FD0EF;
mem['h0F57] = 32'h0E810613;
mem['h0F58] = 32'h08810593;
mem['h0F59] = 32'h10810513;
mem['h0F5A] = 32'hC79FD0EF;
mem['h0F5B] = 32'h0C810613;
mem['h0F5C] = 32'h0A810593;
mem['h0F5D] = 32'h12810513;
mem['h0F5E] = 32'hC69FD0EF;
mem['h0F5F] = 32'h02000613;
mem['h0F60] = 32'h12810593;
mem['h0F61] = 32'h10810513;
mem['h0F62] = 32'hEECFC0EF;
mem['h0F63] = 32'h00051863;
mem['h0F64] = 32'h000065B7;
mem['h0F65] = 32'hC0858593;
mem['h0F66] = 32'hF71FF06F;
mem['h0F67] = 32'h000065B7;
mem['h0F68] = 32'hC5058593;
mem['h0F69] = 32'hF65FF06F;
mem['h0F6A] = 32'h000065B7;
mem['h0F6B] = 32'hC8458593;
mem['h0F6C] = 32'h06810513;
mem['h0F6D] = 32'hF14FC0EF;
mem['h0F6E] = 32'h10051A63;
mem['h0F6F] = 32'h00A00A13;
mem['h0F70] = 32'h00006CB7;
mem['h0F71] = 32'h00005D37;
mem['h0F72] = 32'h02000D93;
mem['h0F73] = 32'h00006B37;
mem['h0F74] = 32'h00006C37;
mem['h0F75] = 32'hC90C8593;
mem['h0F76] = 32'h00040513;
mem['h0F77] = 32'hBE8FC0EF;
mem['h0F78] = 32'h10810513;
mem['h0F79] = 32'hE39FE0EF;
mem['h0F7A] = 32'h01100613;
mem['h0F7B] = 32'h770D0593;
mem['h0F7C] = 32'h12810513;
mem['h0F7D] = 32'h80DFE0EF;
mem['h0F7E] = 32'h00000713;
mem['h0F7F] = 32'h10810793;
mem['h0F80] = 32'h00E787B3;
mem['h0F81] = 32'h0007C783;
mem['h0F82] = 32'h00E12623;
mem['h0F83] = 32'h01010713;
mem['h0F84] = 32'h0047D693;
mem['h0F85] = 32'h00F12423;
mem['h0F86] = 32'h16068793;
mem['h0F87] = 32'h00E786B3;
mem['h0F88] = 32'hFB86C583;
mem['h0F89] = 32'h00040513;
mem['h0F8A] = 32'hA4CFC0EF;
mem['h0F8B] = 32'h00812783;
mem['h0F8C] = 32'h01010713;
mem['h0F8D] = 32'h00040513;
mem['h0F8E] = 32'h00F7F793;
mem['h0F8F] = 32'h16078793;
mem['h0F90] = 32'h00E787B3;
mem['h0F91] = 32'hFB87C583;
mem['h0F92] = 32'hA2CFC0EF;
mem['h0F93] = 32'h00C12703;
mem['h0F94] = 32'h00170713;
mem['h0F95] = 32'hFBB714E3;
mem['h0F96] = 32'hBF0B0593;
mem['h0F97] = 32'h00040513;
mem['h0F98] = 32'hB64FC0EF;
mem['h0F99] = 32'hCB0C0593;
mem['h0F9A] = 32'h00040513;
mem['h0F9B] = 32'hB58FC0EF;
mem['h0F9C] = 32'h12810513;
mem['h0F9D] = 32'hDA9FE0EF;
mem['h0F9E] = 32'h00400613;
mem['h0F9F] = 32'h12810593;
mem['h0FA0] = 32'h0E810513;
mem['h0FA1] = 32'hF7CFE0EF;
mem['h0FA2] = 32'h02000613;
mem['h0FA3] = 32'h00000593;
mem['h0FA4] = 32'h12810513;
mem['h0FA5] = 32'hD88FE0EF;
mem['h0FA6] = 32'h0E812503;
mem['h0FA7] = 32'h3DF00593;
mem['h0FA8] = 32'hFFFA0A13;
mem['h0FA9] = 32'h069010EF;
mem['h0FAA] = 32'h00A50593;
mem['h0FAB] = 32'h00040513;
mem['h0FAC] = 32'hA58FC0EF;
mem['h0FAD] = 32'hBF0B0593;
mem['h0FAE] = 32'h00040513;
mem['h0FAF] = 32'h0FFA7A13;
mem['h0FB0] = 32'hB04FC0EF;
mem['h0FB1] = 32'hF00A18E3;
mem['h0FB2] = 32'hD31FF06F;
mem['h0FB3] = 32'h000065B7;
mem['h0FB4] = 32'hCE058593;
mem['h0FB5] = 32'h06810513;
mem['h0FB6] = 32'hDF0FC0EF;
mem['h0FB7] = 32'h02050463;
mem['h0FB8] = 32'h000065B7;
mem['h0FB9] = 32'hD0458593;
mem['h0FBA] = 32'h06810513;
mem['h0FBB] = 32'hDDCFC0EF;
mem['h0FBC] = 32'h06051263;
mem['h0FBD] = 32'h00040513;
mem['h0FBE] = 32'h8F9FD0EF;
mem['h0FBF] = 32'hCFDFF06F;
mem['h0FC0] = 32'h01C0006F;
mem['h0FC1] = 32'h00014B37;
mem['h0FC2] = 32'h00A00A13;
mem['h0FC3] = 32'h87FB0B13;
mem['h0FC4] = 32'h00006C37;
mem['h0FC5] = 32'h3E800793;
mem['h0FC6] = 32'hC00026F3;
mem['h0FC7] = 32'hC0002773;
mem['h0FC8] = 32'h40D70733;
mem['h0FC9] = 32'hFCEB7EE3;
mem['h0FCA] = 32'hFFF78793;
mem['h0FCB] = 32'hFE0796E3;
mem['h0FCC] = 32'hFFFA0A13;
mem['h0FCD] = 32'hCECC0593;
mem['h0FCE] = 32'h00040513;
mem['h0FCF] = 32'h0FFA7A13;
mem['h0FD0] = 32'hA84FC0EF;
mem['h0FD1] = 32'hFC0A18E3;
mem['h0FD2] = 32'h000065B7;
mem['h0FD3] = 32'hCF058593;
mem['h0FD4] = 32'hDB9FF06F;
mem['h0FD5] = 32'h000065B7;
mem['h0FD6] = 32'hD1458593;
mem['h0FD7] = 32'h06810513;
mem['h0FD8] = 32'hD68FC0EF;
mem['h0FD9] = 32'h18051A63;
mem['h0FDA] = 32'h000065B7;
mem['h0FDB] = 32'hD2458593;
mem['h0FDC] = 32'h00040513;
mem['h0FDD] = 32'hA50FC0EF;
mem['h0FDE] = 32'h000065B7;
mem['h0FDF] = 32'hD4858593;
mem['h0FE0] = 32'h00040513;
mem['h0FE1] = 32'hA40FC0EF;
mem['h0FE2] = 32'h00098593;
mem['h0FE3] = 32'h00040513;
mem['h0FE4] = 32'hA78FC0EF;
mem['h0FE5] = 32'h00006A37;
mem['h0FE6] = 32'h294A0593;
mem['h0FE7] = 32'h00040513;
mem['h0FE8] = 32'hA24FC0EF;
mem['h0FE9] = 32'h12810593;
mem['h0FEA] = 32'h00040513;
mem['h0FEB] = 32'hAD4FC0EF;
mem['h0FEC] = 32'hFE050AE3;
mem['h0FED] = 32'h00098593;
mem['h0FEE] = 32'h12810513;
mem['h0FEF] = 32'hFCDFD0EF;
mem['h0FF0] = 32'h000065B7;
mem['h0FF1] = 32'hD5858593;
mem['h0FF2] = 32'h00040513;
mem['h0FF3] = 32'h9F8FC0EF;
mem['h0FF4] = 32'h00448593;
mem['h0FF5] = 32'h00040513;
mem['h0FF6] = 32'hA30FC0EF;
mem['h0FF7] = 32'h294A0593;
mem['h0FF8] = 32'h00040513;
mem['h0FF9] = 32'h9E0FC0EF;
mem['h0FFA] = 32'h12810593;
mem['h0FFB] = 32'h00040513;
mem['h0FFC] = 32'hA90FC0EF;
mem['h0FFD] = 32'hFE050AE3;
mem['h0FFE] = 32'h80418593;
mem['h0FFF] = 32'h12810513;
mem['h1000] = 32'hF89FD0EF;
mem['h1001] = 32'h000065B7;
mem['h1002] = 32'hD6858593;
mem['h1003] = 32'h00040513;
mem['h1004] = 32'h9B4FC0EF;
mem['h1005] = 32'h12810593;
mem['h1006] = 32'h00040513;
mem['h1007] = 32'hA64FC0EF;
mem['h1008] = 32'hFE050AE3;
mem['h1009] = 32'h12814783;
mem['h100A] = 32'h05900713;
mem['h100B] = 32'h0DF7F793;
mem['h100C] = 32'h00E79A63;
mem['h100D] = 32'h10810513;
mem['h100E] = 32'hBE5FE0EF;
mem['h100F] = 32'h10815783;
mem['h1010] = 32'h00F49623;
mem['h1011] = 32'h000065B7;
mem['h1012] = 32'hD9058593;
mem['h1013] = 32'h00040513;
mem['h1014] = 32'h974FC0EF;
mem['h1015] = 32'h00E48593;
mem['h1016] = 32'h00040513;
mem['h1017] = 32'h9ACFC0EF;
mem['h1018] = 32'h294A0593;
mem['h1019] = 32'h00040513;
mem['h101A] = 32'h95CFC0EF;
mem['h101B] = 32'h12810593;
mem['h101C] = 32'h00040513;
mem['h101D] = 32'hA0CFC0EF;
mem['h101E] = 32'hFE050AE3;
mem['h101F] = 32'h80E18593;
mem['h1020] = 32'h12810513;
mem['h1021] = 32'hF05FD0EF;
mem['h1022] = 32'h000065B7;
mem['h1023] = 32'hDA458593;
mem['h1024] = 32'h00040513;
mem['h1025] = 32'h930FC0EF;
mem['h1026] = 32'h0124C583;
mem['h1027] = 32'h00040513;
mem['h1028] = 32'h868FC0EF;
mem['h1029] = 32'h294A0593;
mem['h102A] = 32'h00040513;
mem['h102B] = 32'h918FC0EF;
mem['h102C] = 32'h12810593;
mem['h102D] = 32'h00040513;
mem['h102E] = 32'h9C8FC0EF;
mem['h102F] = 32'hFE050AE3;
mem['h1030] = 32'h00300693;
mem['h1031] = 32'h00000613;
mem['h1032] = 32'h10810593;
mem['h1033] = 32'h12810513;
mem['h1034] = 32'h10012423;
mem['h1035] = 32'hC28FC0EF;
mem['h1036] = 32'h00050663;
mem['h1037] = 32'h10812783;
mem['h1038] = 32'h00F48923;
mem['h1039] = 32'h000065B7;
mem['h103A] = 32'hDC058593;
mem['h103B] = 32'h00040513;
mem['h103C] = 32'h8D4FC0EF;
mem['h103D] = 32'hE01FF06F;
mem['h103E] = 32'h000065B7;
mem['h103F] = 32'hDE458593;
mem['h1040] = 32'h06810513;
mem['h1041] = 32'hBC4FC0EF;
mem['h1042] = 32'h00050B13;
mem['h1043] = 32'h06051C63;
mem['h1044] = 32'h02442783;
mem['h1045] = 32'h0007A783;
mem['h1046] = 32'h0007A703;
mem['h1047] = 32'h00072783;
mem['h1048] = 32'h0027E793;
mem['h1049] = 32'h00F72023;
mem['h104A] = 32'h02442783;
mem['h104B] = 32'h0007A783;
mem['h104C] = 32'h0007A783;
mem['h104D] = 32'h0007A783;
mem['h104E] = 32'h0017F793;
mem['h104F] = 32'hFE0786E3;
mem['h1050] = 32'h000065B7;
mem['h1051] = 32'hDF458593;
mem['h1052] = 32'h00040513;
mem['h1053] = 32'h878FC0EF;
mem['h1054] = 32'h04000A13;
mem['h1055] = 32'h000B0593;
mem['h1056] = 32'h00040513;
mem['h1057] = 32'h001B0B13;
mem['h1058] = 32'hF89FC0EF;
mem['h1059] = 32'hFF4B18E3;
mem['h105A] = 32'h02442783;
mem['h105B] = 32'h0007A783;
mem['h105C] = 32'h0007A703;
mem['h105D] = 32'h00072783;
mem['h105E] = 32'hFFD7F793;
mem['h105F] = 32'h00F72023;
mem['h1060] = 32'hA79FF06F;
mem['h1061] = 32'h000065B7;
mem['h1062] = 32'hE0858593;
mem['h1063] = 32'h06810513;
mem['h1064] = 32'hB38FC0EF;
mem['h1065] = 32'h34051863;
mem['h1066] = 32'h02442783;
mem['h1067] = 32'h0007A783;
mem['h1068] = 32'h0007A703;
mem['h1069] = 32'h00072783;
mem['h106A] = 32'h0027E793;
mem['h106B] = 32'h00F72023;
mem['h106C] = 32'h02442783;
mem['h106D] = 32'h0007A783;
mem['h106E] = 32'h0007A783;
mem['h106F] = 32'h0007A783;
mem['h1070] = 32'h0017F793;
mem['h1071] = 32'hFE0786E3;
mem['h1072] = 32'h000065B7;
mem['h1073] = 32'hE1858593;
mem['h1074] = 32'h00040513;
mem['h1075] = 32'hFF1FB0EF;
mem['h1076] = 32'h000065B7;
mem['h1077] = 32'hE3C58593;
mem['h1078] = 32'h00040513;
mem['h1079] = 32'hFE1FB0EF;
mem['h107A] = 32'h12810593;
mem['h107B] = 32'h00040513;
mem['h107C] = 32'h890FC0EF;
mem['h107D] = 32'hFE050AE3;
mem['h107E] = 32'h03F00693;
mem['h107F] = 32'h00000613;
mem['h1080] = 32'h08810593;
mem['h1081] = 32'h12810513;
mem['h1082] = 32'h08012423;
mem['h1083] = 32'hAF0FC0EF;
mem['h1084] = 32'h000065B7;
mem['h1085] = 32'hE5858593;
mem['h1086] = 32'h00040513;
mem['h1087] = 32'hFA9FB0EF;
mem['h1088] = 32'h08812C03;
mem['h1089] = 32'h02842783;
mem['h108A] = 32'h0A810593;
mem['h108B] = 32'h002C1A13;
mem['h108C] = 32'h014787B3;
mem['h108D] = 32'h0007A783;
mem['h108E] = 32'h00040513;
mem['h108F] = 32'h00006B37;
mem['h1090] = 32'h0007A783;
mem['h1091] = 32'h0007A683;
mem['h1092] = 32'h0006D783;
mem['h1093] = 32'h00879713;
mem['h1094] = 32'h0087D793;
mem['h1095] = 32'h00F76733;
mem['h1096] = 32'h0006A783;
mem['h1097] = 32'h0AE11523;
mem['h1098] = 32'h0187D693;
mem['h1099] = 32'h0107D793;
mem['h109A] = 32'h0AD10423;
mem['h109B] = 32'h0AF104A3;
mem['h109C] = 32'hF99FB0EF;
mem['h109D] = 32'h294B0593;
mem['h109E] = 32'h00040513;
mem['h109F] = 32'hF49FB0EF;
mem['h10A0] = 32'h12810593;
mem['h10A1] = 32'h00040513;
mem['h10A2] = 32'hFF9FB0EF;
mem['h10A3] = 32'hFE050AE3;
mem['h10A4] = 32'h0A810593;
mem['h10A5] = 32'h12810513;
mem['h10A6] = 32'hCF1FD0EF;
mem['h10A7] = 32'h000065B7;
mem['h10A8] = 32'hD5858593;
mem['h10A9] = 32'h00040513;
mem['h10AA] = 32'hF1DFB0EF;
mem['h10AB] = 32'h02842783;
mem['h10AC] = 32'h0C810593;
mem['h10AD] = 32'h00040513;
mem['h10AE] = 32'h014787B3;
mem['h10AF] = 32'h0007A783;
mem['h10B0] = 32'h0047A783;
mem['h10B1] = 32'h0007A683;
mem['h10B2] = 32'h0006D783;
mem['h10B3] = 32'h00879713;
mem['h10B4] = 32'h0087D793;
mem['h10B5] = 32'h00F76733;
mem['h10B6] = 32'h0006A783;
mem['h10B7] = 32'h0CE11523;
mem['h10B8] = 32'h0187D693;
mem['h10B9] = 32'h0107D793;
mem['h10BA] = 32'h0CD10423;
mem['h10BB] = 32'h0CF104A3;
mem['h10BC] = 32'hF19FB0EF;
mem['h10BD] = 32'h294B0593;
mem['h10BE] = 32'h00040513;
mem['h10BF] = 32'hEC9FB0EF;
mem['h10C0] = 32'h12810593;
mem['h10C1] = 32'h00040513;
mem['h10C2] = 32'hF79FB0EF;
mem['h10C3] = 32'hFE050AE3;
mem['h10C4] = 32'h0C810593;
mem['h10C5] = 32'h12810513;
mem['h10C6] = 32'hC71FD0EF;
mem['h10C7] = 32'h000065B7;
mem['h10C8] = 32'hE7458593;
mem['h10C9] = 32'h00040513;
mem['h10CA] = 32'hE9DFB0EF;
mem['h10CB] = 32'h02842783;
mem['h10CC] = 32'h00040513;
mem['h10CD] = 32'h014787B3;
mem['h10CE] = 32'h0007A783;
mem['h10CF] = 32'h0087A783;
mem['h10D0] = 32'h0007A783;
mem['h10D1] = 32'h0007A583;
mem['h10D2] = 32'h03F5F593;
mem['h10D3] = 32'h0EB12423;
mem['h10D4] = 32'hDB9FB0EF;
mem['h10D5] = 32'h294B0593;
mem['h10D6] = 32'h00040513;
mem['h10D7] = 32'hE69FB0EF;
mem['h10D8] = 32'h12810593;
mem['h10D9] = 32'h00040513;
mem['h10DA] = 32'hF19FB0EF;
mem['h10DB] = 32'hFE050AE3;
mem['h10DC] = 32'h03F00693;
mem['h10DD] = 32'h00000613;
mem['h10DE] = 32'h0E810593;
mem['h10DF] = 32'h12810513;
mem['h10E0] = 32'h97CFC0EF;
mem['h10E1] = 32'h000065B7;
mem['h10E2] = 32'hE8C58593;
mem['h10E3] = 32'h00040513;
mem['h10E4] = 32'hE35FB0EF;
mem['h10E5] = 32'h02842783;
mem['h10E6] = 32'h00040513;
mem['h10E7] = 32'h014787B3;
mem['h10E8] = 32'h0007A783;
mem['h10E9] = 32'h00C7A783;
mem['h10EA] = 32'h0007A783;
mem['h10EB] = 32'h0007A583;
mem['h10EC] = 32'h0075F593;
mem['h10ED] = 32'h10B12423;
mem['h10EE] = 32'hD51FB0EF;
mem['h10EF] = 32'h294B0593;
mem['h10F0] = 32'h00040513;
mem['h10F1] = 32'hE01FB0EF;
mem['h10F2] = 32'h12810593;
mem['h10F3] = 32'h00040513;
mem['h10F4] = 32'hEB1FB0EF;
mem['h10F5] = 32'hFE050AE3;
mem['h10F6] = 32'h10810593;
mem['h10F7] = 32'h00300693;
mem['h10F8] = 32'h00000613;
mem['h10F9] = 32'h12810513;
mem['h10FA] = 32'h914FC0EF;
mem['h10FB] = 32'h0C814783;
mem['h10FC] = 32'h0C914703;
mem['h10FD] = 32'h000065B7;
mem['h10FE] = 32'h01879793;
mem['h10FF] = 32'h01071713;
mem['h1100] = 32'h00E7E7B3;
mem['h1101] = 32'h0CB14703;
mem['h1102] = 32'h00040513;
mem['h1103] = 32'hE9C58593;
mem['h1104] = 32'h00E7E7B3;
mem['h1105] = 32'h0CA14703;
mem['h1106] = 32'h00871713;
mem['h1107] = 32'h00E7E6B3;
mem['h1108] = 32'h02842703;
mem['h1109] = 32'h01470733;
mem['h110A] = 32'h00072783;
mem['h110B] = 32'h0A914703;
mem['h110C] = 32'h0007A783;
mem['h110D] = 32'h01071713;
mem['h110E] = 32'h0007A603;
mem['h110F] = 32'h0A814783;
mem['h1110] = 32'h01879793;
mem['h1111] = 32'h00E7E7B3;
mem['h1112] = 32'h0AB14703;
mem['h1113] = 32'h00E7E7B3;
mem['h1114] = 32'h0AA14703;
mem['h1115] = 32'h00871713;
mem['h1116] = 32'h00E7E7B3;
mem['h1117] = 32'h02842703;
mem['h1118] = 32'h00F62023;
mem['h1119] = 32'h01470733;
mem['h111A] = 32'h00072783;
mem['h111B] = 32'h0E812703;
mem['h111C] = 32'h0047A783;
mem['h111D] = 32'h03F77713;
mem['h111E] = 32'h0007A783;
mem['h111F] = 32'h00D7A023;
mem['h1120] = 32'h02842783;
mem['h1121] = 32'h014787B3;
mem['h1122] = 32'h0007A783;
mem['h1123] = 32'h0087A783;
mem['h1124] = 32'h0007A683;
mem['h1125] = 32'h0006A783;
mem['h1126] = 32'hFC07F793;
mem['h1127] = 32'h00E7E7B3;
mem['h1128] = 32'h00F6A023;
mem['h1129] = 32'h02842783;
mem['h112A] = 32'h10812703;
mem['h112B] = 32'h014787B3;
mem['h112C] = 32'h0007A783;
mem['h112D] = 32'h00777713;
mem['h112E] = 32'h00C7A783;
mem['h112F] = 32'h0007A683;
mem['h1130] = 32'h0006A783;
mem['h1131] = 32'hFF87F793;
mem['h1132] = 32'h00E7E7B3;
mem['h1133] = 32'h00F6A023;
mem['h1134] = 32'hCF5FB0EF;
mem['h1135] = 32'h000C0593;
mem['h1136] = 32'h00040513;
mem['h1137] = 32'hC0DFC0EF;
mem['h1138] = 32'hC89FF06F;
mem['h1139] = 32'h000065B7;
mem['h113A] = 32'hEBC58593;
mem['h113B] = 32'h06810513;
mem['h113C] = 32'hFD9FB0EF;
mem['h113D] = 32'h00050B13;
mem['h113E] = 32'h06051063;
mem['h113F] = 32'h02442783;
mem['h1140] = 32'h0007A783;
mem['h1141] = 32'h0007A703;
mem['h1142] = 32'h00072783;
mem['h1143] = 32'h0027E793;
mem['h1144] = 32'h00F72023;
mem['h1145] = 32'h02442783;
mem['h1146] = 32'h0007A783;
mem['h1147] = 32'h0007A783;
mem['h1148] = 32'h0007A783;
mem['h1149] = 32'h0017F793;
mem['h114A] = 32'hFE0786E3;
mem['h114B] = 32'h000065B7;
mem['h114C] = 32'hED058593;
mem['h114D] = 32'h00040513;
mem['h114E] = 32'hC8DFB0EF;
mem['h114F] = 32'h04000A13;
mem['h1150] = 32'h000B0593;
mem['h1151] = 32'h00040513;
mem['h1152] = 32'h001B0B13;
mem['h1153] = 32'hD19FC0EF;
mem['h1154] = 32'hFF4B18E3;
mem['h1155] = 32'hC15FF06F;
mem['h1156] = 32'h000065B7;
mem['h1157] = 32'hEE458593;
mem['h1158] = 32'h06810513;
mem['h1159] = 32'hF65FB0EF;
mem['h115A] = 32'h00050463;
mem['h115B] = 32'h6DD0006F;
mem['h115C] = 32'h02442783;
mem['h115D] = 32'h0007A783;
mem['h115E] = 32'h0007A703;
mem['h115F] = 32'h00072783;
mem['h1160] = 32'h0027E793;
mem['h1161] = 32'h00F72023;
mem['h1162] = 32'h02442783;
mem['h1163] = 32'h0007A783;
mem['h1164] = 32'h0007A783;
mem['h1165] = 32'h0007A783;
mem['h1166] = 32'h0017F793;
mem['h1167] = 32'hFE0786E3;
mem['h1168] = 32'h000065B7;
mem['h1169] = 32'hEF858593;
mem['h116A] = 32'h00040513;
mem['h116B] = 32'hC19FB0EF;
mem['h116C] = 32'h000065B7;
mem['h116D] = 32'hE3C58593;
mem['h116E] = 32'h00040513;
mem['h116F] = 32'hC09FB0EF;
mem['h1170] = 32'h12810593;
mem['h1171] = 32'h00040513;
mem['h1172] = 32'hCB9FB0EF;
mem['h1173] = 32'hFE050AE3;
mem['h1174] = 32'h03F00693;
mem['h1175] = 32'h00000613;
mem['h1176] = 32'h01010593;
mem['h1177] = 32'h12810513;
mem['h1178] = 32'h00012823;
mem['h1179] = 32'hF19FB0EF;
mem['h117A] = 32'h000065B7;
mem['h117B] = 32'hF1C58593;
mem['h117C] = 32'h00040513;
mem['h117D] = 32'hBD1FB0EF;
mem['h117E] = 32'h01012C83;
mem['h117F] = 32'h02C42783;
mem['h1180] = 32'h00400613;
mem['h1181] = 32'h002C9A13;
mem['h1182] = 32'h014787B3;
mem['h1183] = 32'h0007A783;
mem['h1184] = 32'h00040513;
mem['h1185] = 32'h00006D37;
mem['h1186] = 32'h0007A783;
mem['h1187] = 32'h0007A783;
mem['h1188] = 32'h0007D583;
mem['h1189] = 32'h00B12A23;
mem['h118A] = 32'hA75FB0EF;
mem['h118B] = 32'h02C42783;
mem['h118C] = 32'h00040513;
mem['h118D] = 32'h00800613;
mem['h118E] = 32'h014787B3;
mem['h118F] = 32'h0007A783;
mem['h1190] = 32'h0047A783;
mem['h1191] = 32'h0007A783;
mem['h1192] = 32'h0007A583;
mem['h1193] = 32'h00B12C23;
mem['h1194] = 32'hA4DFB0EF;
mem['h1195] = 32'h294D0593;
mem['h1196] = 32'h00040513;
mem['h1197] = 32'hB69FB0EF;
mem['h1198] = 32'h12810593;
mem['h1199] = 32'h00040513;
mem['h119A] = 32'hC19FB0EF;
mem['h119B] = 32'hFE050AE3;
mem['h119C] = 32'h12810513;
mem['h119D] = 32'hE35FB0EF;
mem['h119E] = 32'h00D00793;
mem['h119F] = 32'h02F51863;
mem['h11A0] = 32'hFFF00613;
mem['h11A1] = 32'h01810593;
mem['h11A2] = 32'h12C10513;
mem['h11A3] = 32'hAC8FD0EF;
mem['h11A4] = 32'h00010637;
mem['h11A5] = 32'h00A00793;
mem['h11A6] = 32'hFFF60613;
mem['h11A7] = 32'h01410593;
mem['h11A8] = 32'h12810513;
mem['h11A9] = 32'h12F10623;
mem['h11AA] = 32'hAACFD0EF;
mem['h11AB] = 32'h000065B7;
mem['h11AC] = 32'hF3458593;
mem['h11AD] = 32'h00040513;
mem['h11AE] = 32'hB0DFB0EF;
mem['h11AF] = 32'h02C42783;
mem['h11B0] = 32'h01C10593;
mem['h11B1] = 32'h00040513;
mem['h11B2] = 32'h014787B3;
mem['h11B3] = 32'h0007A783;
mem['h11B4] = 32'h0087A783;
mem['h11B5] = 32'h0007A683;
mem['h11B6] = 32'h0006D783;
mem['h11B7] = 32'h00879713;
mem['h11B8] = 32'h0087D793;
mem['h11B9] = 32'h00F76733;
mem['h11BA] = 32'h0006A783;
mem['h11BB] = 32'h00E11F23;
mem['h11BC] = 32'h0187D693;
mem['h11BD] = 32'h0107D793;
mem['h11BE] = 32'h00D10E23;
mem['h11BF] = 32'h00F10EA3;
mem['h11C0] = 32'hB09FB0EF;
mem['h11C1] = 32'h294D0593;
mem['h11C2] = 32'h00040513;
mem['h11C3] = 32'hAB9FB0EF;
mem['h11C4] = 32'h12810593;
mem['h11C5] = 32'h00040513;
mem['h11C6] = 32'hB69FB0EF;
mem['h11C7] = 32'hFE050AE3;
mem['h11C8] = 32'h01C10593;
mem['h11C9] = 32'h12810513;
mem['h11CA] = 32'h861FD0EF;
mem['h11CB] = 32'h01D14783;
mem['h11CC] = 32'h01C14C03;
mem['h11CD] = 32'h000065B7;
mem['h11CE] = 32'h01079793;
mem['h11CF] = 32'h018C1C13;
mem['h11D0] = 32'h00FC6C33;
mem['h11D1] = 32'h01F14783;
mem['h11D2] = 32'hF4C58593;
mem['h11D3] = 32'h00040513;
mem['h11D4] = 32'h00FC6C33;
mem['h11D5] = 32'h01E14783;
mem['h11D6] = 32'h00879793;
mem['h11D7] = 32'h00FC6C33;
mem['h11D8] = 32'hA65FB0EF;
mem['h11D9] = 32'h02C42783;
mem['h11DA] = 32'h00040513;
mem['h11DB] = 32'h014787B3;
mem['h11DC] = 32'h0007A783;
mem['h11DD] = 32'h00C7A783;
mem['h11DE] = 32'h0007A783;
mem['h11DF] = 32'h0007D583;
mem['h11E0] = 32'h02B12023;
mem['h11E1] = 32'h985FB0EF;
mem['h11E2] = 32'h294D0593;
mem['h11E3] = 32'h00040513;
mem['h11E4] = 32'hA35FB0EF;
mem['h11E5] = 32'h12810593;
mem['h11E6] = 32'h00040513;
mem['h11E7] = 32'hAE5FB0EF;
mem['h11E8] = 32'hFE050AE3;
mem['h11E9] = 32'h000106B7;
mem['h11EA] = 32'hFFF68693;
mem['h11EB] = 32'h00000613;
mem['h11EC] = 32'h02010593;
mem['h11ED] = 32'h12810513;
mem['h11EE] = 32'hD45FB0EF;
mem['h11EF] = 32'h000065B7;
mem['h11F0] = 32'hF6858593;
mem['h11F1] = 32'h00040513;
mem['h11F2] = 32'h9FDFB0EF;
mem['h11F3] = 32'h02C42783;
mem['h11F4] = 32'h00040513;
mem['h11F5] = 32'h00800613;
mem['h11F6] = 32'h014787B3;
mem['h11F7] = 32'h0007A783;
mem['h11F8] = 32'h0107A783;
mem['h11F9] = 32'h0007A783;
mem['h11FA] = 32'h0007A583;
mem['h11FB] = 32'h02B12223;
mem['h11FC] = 32'h8ADFB0EF;
mem['h11FD] = 32'h294D0593;
mem['h11FE] = 32'h00040513;
mem['h11FF] = 32'h9C9FB0EF;
mem['h1200] = 32'h12810593;
mem['h1201] = 32'h00040513;
mem['h1202] = 32'hA79FB0EF;
mem['h1203] = 32'hFE050AE3;
mem['h1204] = 32'hFFF00613;
mem['h1205] = 32'h02410593;
mem['h1206] = 32'h12810513;
mem['h1207] = 32'h938FD0EF;
mem['h1208] = 32'h000065B7;
mem['h1209] = 32'hF8458593;
mem['h120A] = 32'h00040513;
mem['h120B] = 32'h999FB0EF;
mem['h120C] = 32'h02C42783;
mem['h120D] = 32'h00400613;
mem['h120E] = 32'h00040513;
mem['h120F] = 32'h014787B3;
mem['h1210] = 32'h0007A783;
mem['h1211] = 32'h0147A783;
mem['h1212] = 32'h0007A783;
mem['h1213] = 32'h0007D583;
mem['h1214] = 32'h02B12423;
mem['h1215] = 32'h849FB0EF;
mem['h1216] = 32'h02C42783;
mem['h1217] = 32'h00040513;
mem['h1218] = 32'h00800613;
mem['h1219] = 32'h014787B3;
mem['h121A] = 32'h0007A783;
mem['h121B] = 32'h0187A783;
mem['h121C] = 32'h0007A783;
mem['h121D] = 32'h0007A583;
mem['h121E] = 32'h02B12623;
mem['h121F] = 32'h821FB0EF;
mem['h1220] = 32'h294D0593;
mem['h1221] = 32'h00040513;
mem['h1222] = 32'h93DFB0EF;
mem['h1223] = 32'h12810593;
mem['h1224] = 32'h00040513;
mem['h1225] = 32'h9EDFB0EF;
mem['h1226] = 32'hFE050AE3;
mem['h1227] = 32'h12810513;
mem['h1228] = 32'hC09FB0EF;
mem['h1229] = 32'h00D00793;
mem['h122A] = 32'h02F51863;
mem['h122B] = 32'hFFF00613;
mem['h122C] = 32'h02C10593;
mem['h122D] = 32'h12C10513;
mem['h122E] = 32'h89CFD0EF;
mem['h122F] = 32'h00010637;
mem['h1230] = 32'h00A00793;
mem['h1231] = 32'hFFF60613;
mem['h1232] = 32'h02810593;
mem['h1233] = 32'h12810513;
mem['h1234] = 32'h12F10623;
mem['h1235] = 32'h880FD0EF;
mem['h1236] = 32'h000065B7;
mem['h1237] = 32'hF9C58593;
mem['h1238] = 32'h00040513;
mem['h1239] = 32'h8E1FB0EF;
mem['h123A] = 32'h02C42783;
mem['h123B] = 32'h03010593;
mem['h123C] = 32'h00040513;
mem['h123D] = 32'h014787B3;
mem['h123E] = 32'h0007A783;
mem['h123F] = 32'h01C7A783;
mem['h1240] = 32'h0007A683;
mem['h1241] = 32'h0006D783;
mem['h1242] = 32'h00879713;
mem['h1243] = 32'h0087D793;
mem['h1244] = 32'h00F76733;
mem['h1245] = 32'h0006A783;
mem['h1246] = 32'h02E11923;
mem['h1247] = 32'h0187D693;
mem['h1248] = 32'h0107D793;
mem['h1249] = 32'h02D10823;
mem['h124A] = 32'h02F108A3;
mem['h124B] = 32'h8DDFB0EF;
mem['h124C] = 32'h294D0593;
mem['h124D] = 32'h00040513;
mem['h124E] = 32'h88DFB0EF;
mem['h124F] = 32'h12810593;
mem['h1250] = 32'h00040513;
mem['h1251] = 32'h93DFB0EF;
mem['h1252] = 32'hFE050AE3;
mem['h1253] = 32'h03010593;
mem['h1254] = 32'h12810513;
mem['h1255] = 32'hE34FD0EF;
mem['h1256] = 32'h03114783;
mem['h1257] = 32'h03014B03;
mem['h1258] = 32'h000065B7;
mem['h1259] = 32'h01079793;
mem['h125A] = 32'h018B1B13;
mem['h125B] = 32'h00FB6B33;
mem['h125C] = 32'h03314783;
mem['h125D] = 32'hFB458593;
mem['h125E] = 32'h00040513;
mem['h125F] = 32'h00FB6B33;
mem['h1260] = 32'h03214783;
mem['h1261] = 32'h00879793;
mem['h1262] = 32'h00FB6B33;
mem['h1263] = 32'h839FB0EF;
mem['h1264] = 32'h02C42783;
mem['h1265] = 32'h00040513;
mem['h1266] = 32'h014787B3;
mem['h1267] = 32'h0007A783;
mem['h1268] = 32'h0207A783;
mem['h1269] = 32'h0007A783;
mem['h126A] = 32'h0007D583;
mem['h126B] = 32'h02B12A23;
mem['h126C] = 32'hF58FB0EF;
mem['h126D] = 32'h294D0593;
mem['h126E] = 32'h00040513;
mem['h126F] = 32'h809FB0EF;
mem['h1270] = 32'h12810593;
mem['h1271] = 32'h00040513;
mem['h1272] = 32'h8B9FB0EF;
mem['h1273] = 32'hFE050AE3;
mem['h1274] = 32'h000106B7;
mem['h1275] = 32'hFFF68693;
mem['h1276] = 32'h00000613;
mem['h1277] = 32'h03410593;
mem['h1278] = 32'h12810513;
mem['h1279] = 32'hB19FB0EF;
mem['h127A] = 32'h000065B7;
mem['h127B] = 32'hFD058593;
mem['h127C] = 32'h00040513;
mem['h127D] = 32'hFD0FB0EF;
mem['h127E] = 32'h02C42783;
mem['h127F] = 32'h00040513;
mem['h1280] = 32'h00800613;
mem['h1281] = 32'h014787B3;
mem['h1282] = 32'h0007A783;
mem['h1283] = 32'h0247A783;
mem['h1284] = 32'h0007A783;
mem['h1285] = 32'h0007A583;
mem['h1286] = 32'h02B12C23;
mem['h1287] = 32'hE80FB0EF;
mem['h1288] = 32'h294D0593;
mem['h1289] = 32'h00040513;
mem['h128A] = 32'hF9CFB0EF;
mem['h128B] = 32'h12810593;
mem['h128C] = 32'h00040513;
mem['h128D] = 32'h84DFB0EF;
mem['h128E] = 32'hFE050AE3;
mem['h128F] = 32'hFFF00613;
mem['h1290] = 32'h03810593;
mem['h1291] = 32'h12810513;
mem['h1292] = 32'hF0DFC0EF;
mem['h1293] = 32'h000065B7;
mem['h1294] = 32'hFF058593;
mem['h1295] = 32'h00040513;
mem['h1296] = 32'hF6CFB0EF;
mem['h1297] = 32'h02C42783;
mem['h1298] = 32'h00040513;
mem['h1299] = 32'h00800613;
mem['h129A] = 32'h014787B3;
mem['h129B] = 32'h0007A783;
mem['h129C] = 32'h0287A783;
mem['h129D] = 32'h0007A783;
mem['h129E] = 32'h0007A583;
mem['h129F] = 32'h02B12E23;
mem['h12A0] = 32'hE1CFB0EF;
mem['h12A1] = 32'h294D0593;
mem['h12A2] = 32'h00040513;
mem['h12A3] = 32'hF38FB0EF;
mem['h12A4] = 32'h12810593;
mem['h12A5] = 32'h00040513;
mem['h12A6] = 32'hFE8FB0EF;
mem['h12A7] = 32'hFE050AE3;
mem['h12A8] = 32'hFFF00613;
mem['h12A9] = 32'h03C10593;
mem['h12AA] = 32'h12810513;
mem['h12AB] = 32'hEA9FC0EF;
mem['h12AC] = 32'h000065B7;
mem['h12AD] = 32'h01858593;
mem['h12AE] = 32'h00040513;
mem['h12AF] = 32'hF08FB0EF;
mem['h12B0] = 32'h02C42783;
mem['h12B1] = 32'h00040513;
mem['h12B2] = 32'h00800613;
mem['h12B3] = 32'h014787B3;
mem['h12B4] = 32'h0007A783;
mem['h12B5] = 32'h02C7A783;
mem['h12B6] = 32'h0007A783;
mem['h12B7] = 32'h0007A583;
mem['h12B8] = 32'h04B12023;
mem['h12B9] = 32'hDB8FB0EF;
mem['h12BA] = 32'h294D0593;
mem['h12BB] = 32'h00040513;
mem['h12BC] = 32'hED4FB0EF;
mem['h12BD] = 32'h12810593;
mem['h12BE] = 32'h00040513;
mem['h12BF] = 32'hF84FB0EF;
mem['h12C0] = 32'hFE050AE3;
mem['h12C1] = 32'hFFF00613;
mem['h12C2] = 32'h04010593;
mem['h12C3] = 32'h12810513;
mem['h12C4] = 32'hE45FC0EF;
mem['h12C5] = 32'h000065B7;
mem['h12C6] = 32'h04058593;
mem['h12C7] = 32'h00040513;
mem['h12C8] = 32'hEA4FB0EF;
mem['h12C9] = 32'h02C42783;
mem['h12CA] = 32'h00040513;
mem['h12CB] = 32'h00800613;
mem['h12CC] = 32'h014787B3;
mem['h12CD] = 32'h0007A783;
mem['h12CE] = 32'h0307A783;
mem['h12CF] = 32'h0007A783;
mem['h12D0] = 32'h0007A583;
mem['h12D1] = 32'h04B12223;
mem['h12D2] = 32'hD54FB0EF;
mem['h12D3] = 32'h294D0593;
mem['h12D4] = 32'h00040513;
mem['h12D5] = 32'hE70FB0EF;
mem['h12D6] = 32'h12810593;
mem['h12D7] = 32'h00040513;
mem['h12D8] = 32'hF20FB0EF;
mem['h12D9] = 32'hFE050AE3;
mem['h12DA] = 32'hFFF00613;
mem['h12DB] = 32'h04410593;
mem['h12DC] = 32'h12810513;
mem['h12DD] = 32'hDE1FC0EF;
mem['h12DE] = 32'h000065B7;
mem['h12DF] = 32'h06858593;
mem['h12E0] = 32'h00040513;
mem['h12E1] = 32'hE40FB0EF;
mem['h12E2] = 32'h02C42783;
mem['h12E3] = 32'h00040513;
mem['h12E4] = 32'h00800613;
mem['h12E5] = 32'h014787B3;
mem['h12E6] = 32'h0007A783;
mem['h12E7] = 32'h0347A783;
mem['h12E8] = 32'h0007A783;
mem['h12E9] = 32'h0007A583;
mem['h12EA] = 32'h04B12423;
mem['h12EB] = 32'hCF0FB0EF;
mem['h12EC] = 32'h294D0593;
mem['h12ED] = 32'h00040513;
mem['h12EE] = 32'hE0CFB0EF;
mem['h12EF] = 32'h12810593;
mem['h12F0] = 32'h00040513;
mem['h12F1] = 32'hEBCFB0EF;
mem['h12F2] = 32'hFE050AE3;
mem['h12F3] = 32'hFFF00613;
mem['h12F4] = 32'h04810593;
mem['h12F5] = 32'h12810513;
mem['h12F6] = 32'hD7DFC0EF;
mem['h12F7] = 32'h000065B7;
mem['h12F8] = 32'h09058593;
mem['h12F9] = 32'h00040513;
mem['h12FA] = 32'hDDCFB0EF;
mem['h12FB] = 32'h02C42783;
mem['h12FC] = 32'h00040513;
mem['h12FD] = 32'h00800613;
mem['h12FE] = 32'h014787B3;
mem['h12FF] = 32'h0007A783;
mem['h1300] = 32'h0387A783;
mem['h1301] = 32'h0007A783;
mem['h1302] = 32'h0007A583;
mem['h1303] = 32'h04B12623;
mem['h1304] = 32'hC8CFB0EF;
mem['h1305] = 32'h294D0593;
mem['h1306] = 32'h00040513;
mem['h1307] = 32'hDA8FB0EF;
mem['h1308] = 32'h12810593;
mem['h1309] = 32'h00040513;
mem['h130A] = 32'hE58FB0EF;
mem['h130B] = 32'hFE050AE3;
mem['h130C] = 32'hFFF00613;
mem['h130D] = 32'h04C10593;
mem['h130E] = 32'h12810513;
mem['h130F] = 32'hD19FC0EF;
mem['h1310] = 32'h000065B7;
mem['h1311] = 32'h0B858593;
mem['h1312] = 32'h00040513;
mem['h1313] = 32'hD78FB0EF;
mem['h1314] = 32'h02C42783;
mem['h1315] = 32'h00040513;
mem['h1316] = 32'h00800613;
mem['h1317] = 32'h014787B3;
mem['h1318] = 32'h0007A783;
mem['h1319] = 32'h03C7A783;
mem['h131A] = 32'h0007A783;
mem['h131B] = 32'h0007A583;
mem['h131C] = 32'h04B12823;
mem['h131D] = 32'hC28FB0EF;
mem['h131E] = 32'h294D0593;
mem['h131F] = 32'h00040513;
mem['h1320] = 32'hD44FB0EF;
mem['h1321] = 32'h12810593;
mem['h1322] = 32'h00040513;
mem['h1323] = 32'hDF4FB0EF;
mem['h1324] = 32'hFE050AE3;
mem['h1325] = 32'hFFF00613;
mem['h1326] = 32'h05010593;
mem['h1327] = 32'h12810513;
mem['h1328] = 32'hCB5FC0EF;
mem['h1329] = 32'h000065B7;
mem['h132A] = 32'h0E058593;
mem['h132B] = 32'h00040513;
mem['h132C] = 32'hD14FB0EF;
mem['h132D] = 32'h02C42783;
mem['h132E] = 32'h00040513;
mem['h132F] = 32'h00800613;
mem['h1330] = 32'h014787B3;
mem['h1331] = 32'h0007A783;
mem['h1332] = 32'h0407A783;
mem['h1333] = 32'h0007A783;
mem['h1334] = 32'h0007A583;
mem['h1335] = 32'h04B12A23;
mem['h1336] = 32'hBC4FB0EF;
mem['h1337] = 32'h294D0593;
mem['h1338] = 32'h00040513;
mem['h1339] = 32'hCE0FB0EF;
mem['h133A] = 32'h12810593;
mem['h133B] = 32'h00040513;
mem['h133C] = 32'hD90FB0EF;
mem['h133D] = 32'hFE050AE3;
mem['h133E] = 32'hFFF00613;
mem['h133F] = 32'h05410593;
mem['h1340] = 32'h12810513;
mem['h1341] = 32'hC51FC0EF;
mem['h1342] = 32'h000065B7;
mem['h1343] = 32'h10858593;
mem['h1344] = 32'h00040513;
mem['h1345] = 32'hCB0FB0EF;
mem['h1346] = 32'h02C42783;
mem['h1347] = 32'h002C9A13;
mem['h1348] = 32'h00040513;
mem['h1349] = 32'h014787B3;
mem['h134A] = 32'h0007A783;
mem['h134B] = 32'h00800613;
mem['h134C] = 32'h00006D37;
mem['h134D] = 32'h0447A783;
mem['h134E] = 32'h0007A783;
mem['h134F] = 32'h0007A583;
mem['h1350] = 32'h04B12C23;
mem['h1351] = 32'hB58FB0EF;
mem['h1352] = 32'h294D0593;
mem['h1353] = 32'h00040513;
mem['h1354] = 32'hC74FB0EF;
mem['h1355] = 32'h12810593;
mem['h1356] = 32'h00040513;
mem['h1357] = 32'hD24FB0EF;
mem['h1358] = 32'hFE050AE3;
mem['h1359] = 32'hFFF00613;
mem['h135A] = 32'h05810593;
mem['h135B] = 32'h12810513;
mem['h135C] = 32'hBE5FC0EF;
mem['h135D] = 32'h000065B7;
mem['h135E] = 32'h13058593;
mem['h135F] = 32'h00040513;
mem['h1360] = 32'hC44FB0EF;
mem['h1361] = 32'h02C42783;
mem['h1362] = 32'h00040513;
mem['h1363] = 32'h00800613;
mem['h1364] = 32'h014787B3;
mem['h1365] = 32'h0007A783;
mem['h1366] = 32'h0487A783;
mem['h1367] = 32'h0007A783;
mem['h1368] = 32'h0007A583;
mem['h1369] = 32'h04B12E23;
mem['h136A] = 32'hAF4FB0EF;
mem['h136B] = 32'h294D0593;
mem['h136C] = 32'h00040513;
mem['h136D] = 32'hC10FB0EF;
mem['h136E] = 32'h12810593;
mem['h136F] = 32'h00040513;
mem['h1370] = 32'hCC0FB0EF;
mem['h1371] = 32'hFE050AE3;
mem['h1372] = 32'hFFF00613;
mem['h1373] = 32'h05C10593;
mem['h1374] = 32'h12810513;
mem['h1375] = 32'hB81FC0EF;
mem['h1376] = 32'h000065B7;
mem['h1377] = 32'h15858593;
mem['h1378] = 32'h00040513;
mem['h1379] = 32'hBE0FB0EF;
mem['h137A] = 32'h02C42783;
mem['h137B] = 32'h00040513;
mem['h137C] = 32'h00800613;
mem['h137D] = 32'h014787B3;
mem['h137E] = 32'h0007A783;
mem['h137F] = 32'h04C7A783;
mem['h1380] = 32'h0007A783;
mem['h1381] = 32'h0007A583;
mem['h1382] = 32'h06B12023;
mem['h1383] = 32'hA90FB0EF;
mem['h1384] = 32'h294D0593;
mem['h1385] = 32'h00040513;
mem['h1386] = 32'hBACFB0EF;
mem['h1387] = 32'h12810593;
mem['h1388] = 32'h00040513;
mem['h1389] = 32'hC5CFB0EF;
mem['h138A] = 32'hFE050AE3;
mem['h138B] = 32'hFFF00613;
mem['h138C] = 32'h06010593;
mem['h138D] = 32'h12810513;
mem['h138E] = 32'hB1DFC0EF;
mem['h138F] = 32'h000065B7;
mem['h1390] = 32'h18058593;
mem['h1391] = 32'h00040513;
mem['h1392] = 32'hB7CFB0EF;
mem['h1393] = 32'h02C42783;
mem['h1394] = 32'h00040513;
mem['h1395] = 32'h00800613;
mem['h1396] = 32'h014787B3;
mem['h1397] = 32'h0007A783;
mem['h1398] = 32'h0507A783;
mem['h1399] = 32'h0007A783;
mem['h139A] = 32'h0007A583;
mem['h139B] = 32'h06B12223;
mem['h139C] = 32'hA2CFB0EF;
mem['h139D] = 32'h294D0593;
mem['h139E] = 32'h00040513;
mem['h139F] = 32'hB48FB0EF;
mem['h13A0] = 32'h12810593;
mem['h13A1] = 32'h00040513;
mem['h13A2] = 32'hBF8FB0EF;
mem['h13A3] = 32'hFE050AE3;
mem['h13A4] = 32'hFFF00613;
mem['h13A5] = 32'h06410593;
mem['h13A6] = 32'h12810513;
mem['h13A7] = 32'hAB9FC0EF;
mem['h13A8] = 32'h000065B7;
mem['h13A9] = 32'h1A858593;
mem['h13AA] = 32'h00040513;
mem['h13AB] = 32'hB18FB0EF;
mem['h13AC] = 32'h02C42783;
mem['h13AD] = 32'h00040513;
mem['h13AE] = 32'h00800613;
mem['h13AF] = 32'h014787B3;
mem['h13B0] = 32'h0007A783;
mem['h13B1] = 32'h0547A783;
mem['h13B2] = 32'h0007A783;
mem['h13B3] = 32'h0007A583;
mem['h13B4] = 32'h08B12423;
mem['h13B5] = 32'h9C8FB0EF;
mem['h13B6] = 32'h294D0593;
mem['h13B7] = 32'h00040513;
mem['h13B8] = 32'hAE4FB0EF;
mem['h13B9] = 32'h12810593;
mem['h13BA] = 32'h00040513;
mem['h13BB] = 32'hB94FB0EF;
mem['h13BC] = 32'hFE050AE3;
mem['h13BD] = 32'hFFF00613;
mem['h13BE] = 32'h08810593;
mem['h13BF] = 32'h12810513;
mem['h13C0] = 32'hA55FC0EF;
mem['h13C1] = 32'h000065B7;
mem['h13C2] = 32'h1D058593;
mem['h13C3] = 32'h00040513;
mem['h13C4] = 32'hAB4FB0EF;
mem['h13C5] = 32'h02C42783;
mem['h13C6] = 32'h00040513;
mem['h13C7] = 32'h00800613;
mem['h13C8] = 32'h014787B3;
mem['h13C9] = 32'h0007A783;
mem['h13CA] = 32'h0587A783;
mem['h13CB] = 32'h0007A783;
mem['h13CC] = 32'h0007A583;
mem['h13CD] = 32'h0AB12423;
mem['h13CE] = 32'h964FB0EF;
mem['h13CF] = 32'h294D0593;
mem['h13D0] = 32'h00040513;
mem['h13D1] = 32'hA80FB0EF;
mem['h13D2] = 32'h12810593;
mem['h13D3] = 32'h00040513;
mem['h13D4] = 32'hB30FB0EF;
mem['h13D5] = 32'hFE050AE3;
mem['h13D6] = 32'hFFF00613;
mem['h13D7] = 32'h0A810593;
mem['h13D8] = 32'h12810513;
mem['h13D9] = 32'h9F1FC0EF;
mem['h13DA] = 32'h000065B7;
mem['h13DB] = 32'h1F858593;
mem['h13DC] = 32'h00040513;
mem['h13DD] = 32'hA50FB0EF;
mem['h13DE] = 32'h02C42783;
mem['h13DF] = 32'h00040513;
mem['h13E0] = 32'h00800613;
mem['h13E1] = 32'h014787B3;
mem['h13E2] = 32'h0007A783;
mem['h13E3] = 32'h05C7A783;
mem['h13E4] = 32'h0007A783;
mem['h13E5] = 32'h0007A583;
mem['h13E6] = 32'h0CB12423;
mem['h13E7] = 32'h900FB0EF;
mem['h13E8] = 32'h294D0593;
mem['h13E9] = 32'h00040513;
mem['h13EA] = 32'hA1CFB0EF;
mem['h13EB] = 32'h12810593;
mem['h13EC] = 32'h00040513;
mem['h13ED] = 32'hACCFB0EF;
mem['h13EE] = 32'hFE050AE3;
mem['h13EF] = 32'hFFF00613;
mem['h13F0] = 32'h0C810593;
mem['h13F1] = 32'h12810513;
mem['h13F2] = 32'h98DFC0EF;
mem['h13F3] = 32'h000065B7;
mem['h13F4] = 32'h22058593;
mem['h13F5] = 32'h00040513;
mem['h13F6] = 32'h9ECFB0EF;
mem['h13F7] = 32'h02C42783;
mem['h13F8] = 32'h00040513;
mem['h13F9] = 32'h00800613;
mem['h13FA] = 32'h014787B3;
mem['h13FB] = 32'h0007A783;
mem['h13FC] = 32'h0607A783;
mem['h13FD] = 32'h0007A783;
mem['h13FE] = 32'h0007A583;
mem['h13FF] = 32'h0EB12423;
mem['h1400] = 32'h89CFB0EF;
mem['h1401] = 32'h294D0593;
mem['h1402] = 32'h00040513;
mem['h1403] = 32'h9B8FB0EF;
mem['h1404] = 32'h12810593;
mem['h1405] = 32'h00040513;
mem['h1406] = 32'hA68FB0EF;
mem['h1407] = 32'hFE050AE3;
mem['h1408] = 32'hFFF00613;
mem['h1409] = 32'h0E810593;
mem['h140A] = 32'h12810513;
mem['h140B] = 32'h929FC0EF;
mem['h140C] = 32'h000065B7;
mem['h140D] = 32'h24858593;
mem['h140E] = 32'h00040513;
mem['h140F] = 32'h988FB0EF;
mem['h1410] = 32'h02C42783;
mem['h1411] = 32'h00040513;
mem['h1412] = 32'h00800613;
mem['h1413] = 32'h014787B3;
mem['h1414] = 32'h0007A783;
mem['h1415] = 32'h0647A783;
mem['h1416] = 32'h0007A783;
mem['h1417] = 32'h0007A583;
mem['h1418] = 32'h10B12423;
mem['h1419] = 32'h838FB0EF;
mem['h141A] = 32'h294D0593;
mem['h141B] = 32'h00040513;
mem['h141C] = 32'h954FB0EF;
mem['h141D] = 32'h12810593;
mem['h141E] = 32'h00040513;
mem['h141F] = 32'hA04FB0EF;
mem['h1420] = 32'hFE050AE3;
mem['h1421] = 32'hFFF00613;
mem['h1422] = 32'h10810593;
mem['h1423] = 32'h12810513;
mem['h1424] = 32'h8C5FC0EF;
mem['h1425] = 32'h02C42783;
mem['h1426] = 32'h01415603;
mem['h1427] = 32'hFFFF0737;
mem['h1428] = 32'h014787B3;
mem['h1429] = 32'h0007A783;
mem['h142A] = 32'h000065B7;
mem['h142B] = 32'h27058593;
mem['h142C] = 32'h0007A783;
mem['h142D] = 32'h00040513;
mem['h142E] = 32'h0007A683;
mem['h142F] = 32'h0006A783;
mem['h1430] = 32'h00E7F7B3;
mem['h1431] = 32'h00C7E7B3;
mem['h1432] = 32'h00F6A023;
mem['h1433] = 32'h02C42783;
mem['h1434] = 32'h01812683;
mem['h1435] = 32'h02015603;
mem['h1436] = 32'h014787B3;
mem['h1437] = 32'h0007A783;
mem['h1438] = 32'h0047A783;
mem['h1439] = 32'h0007A783;
mem['h143A] = 32'h00D7A023;
mem['h143B] = 32'h02C42783;
mem['h143C] = 32'h014787B3;
mem['h143D] = 32'h0007A783;
mem['h143E] = 32'h0087A783;
mem['h143F] = 32'h0007A783;
mem['h1440] = 32'h0187A023;
mem['h1441] = 32'h02C42783;
mem['h1442] = 32'h014787B3;
mem['h1443] = 32'h0007A783;
mem['h1444] = 32'h00C7A783;
mem['h1445] = 32'h0007A683;
mem['h1446] = 32'h0006A783;
mem['h1447] = 32'h00E7F7B3;
mem['h1448] = 32'h00C7E7B3;
mem['h1449] = 32'h00F6A023;
mem['h144A] = 32'h02C42783;
mem['h144B] = 32'h02412683;
mem['h144C] = 32'h014787B3;
mem['h144D] = 32'h0007A783;
mem['h144E] = 32'h0107A783;
mem['h144F] = 32'h0007A783;
mem['h1450] = 32'h00D7A023;
mem['h1451] = 32'h02C42783;
mem['h1452] = 32'h014787B3;
mem['h1453] = 32'h0007A783;
mem['h1454] = 32'h02815603;
mem['h1455] = 32'h0147A783;
mem['h1456] = 32'h0007A683;
mem['h1457] = 32'h0006A783;
mem['h1458] = 32'h00E7F7B3;
mem['h1459] = 32'h00C7E7B3;
mem['h145A] = 32'h00F6A023;
mem['h145B] = 32'h02C42783;
mem['h145C] = 32'h02C12683;
mem['h145D] = 32'h03415603;
mem['h145E] = 32'h014787B3;
mem['h145F] = 32'h0007A783;
mem['h1460] = 32'h0187A783;
mem['h1461] = 32'h0007A783;
mem['h1462] = 32'h00D7A023;
mem['h1463] = 32'h02C42783;
mem['h1464] = 32'h014787B3;
mem['h1465] = 32'h0007A783;
mem['h1466] = 32'h01C7A783;
mem['h1467] = 32'h0007A783;
mem['h1468] = 32'h0167A023;
mem['h1469] = 32'h02C42783;
mem['h146A] = 32'h014787B3;
mem['h146B] = 32'h0007A783;
mem['h146C] = 32'h0207A783;
mem['h146D] = 32'h0007A683;
mem['h146E] = 32'h0006A783;
mem['h146F] = 32'h00E7F7B3;
mem['h1470] = 32'h00C7E7B3;
mem['h1471] = 32'h00F6A023;
mem['h1472] = 32'h02C42783;
mem['h1473] = 32'h03812703;
mem['h1474] = 32'h014787B3;
mem['h1475] = 32'h0007A783;
mem['h1476] = 32'h0247A783;
mem['h1477] = 32'h0007A783;
mem['h1478] = 32'h00E7A023;
mem['h1479] = 32'h02C42783;
mem['h147A] = 32'h014787B3;
mem['h147B] = 32'h0007A783;
mem['h147C] = 32'h0287A783;
mem['h147D] = 32'h03C12703;
mem['h147E] = 32'h0007A783;
mem['h147F] = 32'h00E7A023;
mem['h1480] = 32'h02C42783;
mem['h1481] = 32'h04012703;
mem['h1482] = 32'h014787B3;
mem['h1483] = 32'h0007A783;
mem['h1484] = 32'h02C7A783;
mem['h1485] = 32'h0007A783;
mem['h1486] = 32'h00E7A023;
mem['h1487] = 32'h02C42783;
mem['h1488] = 32'h04412703;
mem['h1489] = 32'h014787B3;
mem['h148A] = 32'h0007A783;
mem['h148B] = 32'h0307A783;
mem['h148C] = 32'h0007A783;
mem['h148D] = 32'h00E7A023;
mem['h148E] = 32'h02C42783;
mem['h148F] = 32'h04812703;
mem['h1490] = 32'h014787B3;
mem['h1491] = 32'h0007A783;
mem['h1492] = 32'h0347A783;
mem['h1493] = 32'h0007A783;
mem['h1494] = 32'h00E7A023;
mem['h1495] = 32'h02C42783;
mem['h1496] = 32'h04C12703;
mem['h1497] = 32'h014787B3;
mem['h1498] = 32'h0007A783;
mem['h1499] = 32'h0387A783;
mem['h149A] = 32'h0007A783;
mem['h149B] = 32'h00E7A023;
mem['h149C] = 32'h02C42783;
mem['h149D] = 32'h014787B3;
mem['h149E] = 32'h0007A783;
mem['h149F] = 32'h03C7A783;
mem['h14A0] = 32'h0007A783;
mem['h14A1] = 32'h05012703;
mem['h14A2] = 32'h00E7A023;
mem['h14A3] = 32'h02C42783;
mem['h14A4] = 32'h05412703;
mem['h14A5] = 32'h014787B3;
mem['h14A6] = 32'h0007A783;
mem['h14A7] = 32'h0407A783;
mem['h14A8] = 32'h0007A783;
mem['h14A9] = 32'h00E7A023;
mem['h14AA] = 32'h02C42783;
mem['h14AB] = 32'h05812703;
mem['h14AC] = 32'h014787B3;
mem['h14AD] = 32'h0007A783;
mem['h14AE] = 32'h0447A783;
mem['h14AF] = 32'h0007A783;
mem['h14B0] = 32'h00E7A023;
mem['h14B1] = 32'h02C42783;
mem['h14B2] = 32'h05C12703;
mem['h14B3] = 32'h014787B3;
mem['h14B4] = 32'h0007A783;
mem['h14B5] = 32'h0487A783;
mem['h14B6] = 32'h0007A783;
mem['h14B7] = 32'h00E7A023;
mem['h14B8] = 32'h02C42783;
mem['h14B9] = 32'h06012703;
mem['h14BA] = 32'h014787B3;
mem['h14BB] = 32'h0007A783;
mem['h14BC] = 32'h04C7A783;
mem['h14BD] = 32'h0007A783;
mem['h14BE] = 32'h00E7A023;
mem['h14BF] = 32'h02C42783;
mem['h14C0] = 32'h06412703;
mem['h14C1] = 32'h014787B3;
mem['h14C2] = 32'h0007A783;
mem['h14C3] = 32'h0507A783;
mem['h14C4] = 32'h0007A783;
mem['h14C5] = 32'h00E7A023;
mem['h14C6] = 32'h02C42783;
mem['h14C7] = 32'h08812703;
mem['h14C8] = 32'h014787B3;
mem['h14C9] = 32'h0007A783;
mem['h14CA] = 32'h0547A783;
mem['h14CB] = 32'h0007A783;
mem['h14CC] = 32'h00E7A023;
mem['h14CD] = 32'h02C42783;
mem['h14CE] = 32'h0A812703;
mem['h14CF] = 32'h014787B3;
mem['h14D0] = 32'h0007A783;
mem['h14D1] = 32'h0587A783;
mem['h14D2] = 32'h0007A783;
mem['h14D3] = 32'h00E7A023;
mem['h14D4] = 32'h02C42783;
mem['h14D5] = 32'h0C812703;
mem['h14D6] = 32'h014787B3;
mem['h14D7] = 32'h0007A783;
mem['h14D8] = 32'h05C7A783;
mem['h14D9] = 32'h0007A783;
mem['h14DA] = 32'h00E7A023;
mem['h14DB] = 32'h02C42783;
mem['h14DC] = 32'h0E812703;
mem['h14DD] = 32'h014787B3;
mem['h14DE] = 32'h0007A783;
mem['h14DF] = 32'h0607A783;
mem['h14E0] = 32'h0007A783;
mem['h14E1] = 32'h00E7A023;
mem['h14E2] = 32'h02C42783;
mem['h14E3] = 32'h10812703;
mem['h14E4] = 32'h014787B3;
mem['h14E5] = 32'h0007A783;
mem['h14E6] = 32'h0647A783;
mem['h14E7] = 32'h0007A783;
mem['h14E8] = 32'h00E7A023;
mem['h14E9] = 32'hE21FA0EF;
mem['h14EA] = 32'h12810593;
mem['h14EB] = 32'h00040513;
mem['h14EC] = 32'hED1FA0EF;
mem['h14ED] = 32'hFE050AE3;
mem['h14EE] = 32'h12814783;
mem['h14EF] = 32'h05900713;
mem['h14F0] = 32'h0DF7F793;
mem['h14F1] = 32'h06E79263;
mem['h14F2] = 32'h02C42783;
mem['h14F3] = 32'h014787B3;
mem['h14F4] = 32'h0007A783;
mem['h14F5] = 32'h0687A783;
mem['h14F6] = 32'h0007A783;
mem['h14F7] = 32'h0007A023;
mem['h14F8] = 32'h02C42783;
mem['h14F9] = 32'h014787B3;
mem['h14FA] = 32'h0007A783;
mem['h14FB] = 32'h06C7A783;
mem['h14FC] = 32'h0007A783;
mem['h14FD] = 32'h0007A023;
mem['h14FE] = 32'h02C42783;
mem['h14FF] = 32'h014787B3;
mem['h1500] = 32'h0007A783;
mem['h1501] = 32'h0707A783;
mem['h1502] = 32'h0007A783;
mem['h1503] = 32'h0007A023;
mem['h1504] = 32'h02C42783;
mem['h1505] = 32'h014787B3;
mem['h1506] = 32'h0007A783;
mem['h1507] = 32'h0747A783;
mem['h1508] = 32'h0007A783;
mem['h1509] = 32'h0007A023;
mem['h150A] = 32'h000065B7;
mem['h150B] = 32'h00040513;
mem['h150C] = 32'h29858593;
mem['h150D] = 32'hD91FA0EF;
mem['h150E] = 32'h000C8593;
mem['h150F] = 32'h00040513;
mem['h1510] = 32'hE25FB0EF;
mem['h1511] = 32'hD25FE06F;
mem['h1512] = 32'h000065B7;
mem['h1513] = 32'h2BC58593;
mem['h1514] = 32'h06810513;
mem['h1515] = 32'h874FB0EF;
mem['h1516] = 32'h04051463;
mem['h1517] = 32'h000065B7;
mem['h1518] = 32'h2C458593;
mem['h1519] = 32'h00040513;
mem['h151A] = 32'hD5DFA0EF;
mem['h151B] = 32'h00091E63;
mem['h151C] = 32'h000065B7;
mem['h151D] = 32'h2D058593;
mem['h151E] = 32'h00040513;
mem['h151F] = 32'hD49FA0EF;
mem['h1520] = 32'h00100913;
mem['h1521] = 32'hF74FE06F;
mem['h1522] = 32'h000065B7;
mem['h1523] = 32'h2DC58593;
mem['h1524] = 32'h00040513;
mem['h1525] = 32'hD31FA0EF;
mem['h1526] = 32'h00000913;
mem['h1527] = 32'hF5CFE06F;
mem['h1528] = 32'h000065B7;
mem['h1529] = 32'h2E858593;
mem['h152A] = 32'h06810513;
mem['h152B] = 32'h81CFB0EF;
mem['h152C] = 32'h00051663;
mem['h152D] = 32'h00000067;
mem['h152E] = 32'hF40FE06F;
mem['h152F] = 32'h000065B7;
mem['h1530] = 32'h2F058593;
mem['h1531] = 32'h06810513;
mem['h1532] = 32'h800FB0EF;
mem['h1533] = 32'h0E051863;
mem['h1534] = 32'h000065B7;
mem['h1535] = 32'h2F858593;
mem['h1536] = 32'h00040513;
mem['h1537] = 32'hCE9FA0EF;
mem['h1538] = 32'h000065B7;
mem['h1539] = 32'h31058593;
mem['h153A] = 32'h00040513;
mem['h153B] = 32'hCD9FA0EF;
mem['h153C] = 32'h000065B7;
mem['h153D] = 32'h34C58593;
mem['h153E] = 32'h00040513;
mem['h153F] = 32'hCC9FA0EF;
mem['h1540] = 32'h000065B7;
mem['h1541] = 32'h38458593;
mem['h1542] = 32'h00040513;
mem['h1543] = 32'hCB9FA0EF;
mem['h1544] = 32'h000065B7;
mem['h1545] = 32'h3C058593;
mem['h1546] = 32'h00040513;
mem['h1547] = 32'hCA9FA0EF;
mem['h1548] = 32'h000065B7;
mem['h1549] = 32'h3FC58593;
mem['h154A] = 32'h00040513;
mem['h154B] = 32'hC99FA0EF;
mem['h154C] = 32'h000065B7;
mem['h154D] = 32'h43458593;
mem['h154E] = 32'h00040513;
mem['h154F] = 32'hC89FA0EF;
mem['h1550] = 32'h000065B7;
mem['h1551] = 32'h46C58593;
mem['h1552] = 32'h00040513;
mem['h1553] = 32'hC79FA0EF;
mem['h1554] = 32'h000065B7;
mem['h1555] = 32'h4A458593;
mem['h1556] = 32'h00040513;
mem['h1557] = 32'hC69FA0EF;
mem['h1558] = 32'h000065B7;
mem['h1559] = 32'h4D458593;
mem['h155A] = 32'h00040513;
mem['h155B] = 32'hC59FA0EF;
mem['h155C] = 32'h000065B7;
mem['h155D] = 32'h51058593;
mem['h155E] = 32'h00040513;
mem['h155F] = 32'hC49FA0EF;
mem['h1560] = 32'h000065B7;
mem['h1561] = 32'h54458593;
mem['h1562] = 32'h00040513;
mem['h1563] = 32'hC39FA0EF;
mem['h1564] = 32'h000065B7;
mem['h1565] = 32'h58458593;
mem['h1566] = 32'h00040513;
mem['h1567] = 32'hC29FA0EF;
mem['h1568] = 32'h000065B7;
mem['h1569] = 32'h5B458593;
mem['h156A] = 32'h00040513;
mem['h156B] = 32'hC19FA0EF;
mem['h156C] = 32'h000065B7;
mem['h156D] = 32'h5E458593;
mem['h156E] = 32'hF50FE06F;
mem['h156F] = 32'h00100793;
mem['h1570] = 32'h00FA1463;
mem['h1571] = 32'hE34FE06F;
mem['h1572] = 32'h000065B7;
mem['h1573] = 32'h61858593;
mem['h1574] = 32'hF38FE06F;
mem['h1575] = 32'h02060063;
mem['h1576] = 32'h02000793;
mem['h1577] = 32'h40C787B3;
mem['h1578] = 32'h00F04C63;
mem['h1579] = 32'hFE060613;
mem['h157A] = 32'h00C515B3;
mem['h157B] = 32'h00000713;
mem['h157C] = 32'h00070513;
mem['h157D] = 32'h00008067;
mem['h157E] = 32'h00C51733;
mem['h157F] = 32'h00C595B3;
mem['h1580] = 32'h00F55533;
mem['h1581] = 32'h00A5E5B3;
mem['h1582] = 32'hFE9FF06F;
mem['h1583] = 32'h00050613;
mem['h1584] = 32'h00000513;
mem['h1585] = 32'h0015F693;
mem['h1586] = 32'h00068463;
mem['h1587] = 32'h00C50533;
mem['h1588] = 32'h0015D593;
mem['h1589] = 32'h00161613;
mem['h158A] = 32'hFE0596E3;
mem['h158B] = 32'h00008067;
mem['h158C] = 32'h00050E13;
mem['h158D] = 32'hFF010113;
mem['h158E] = 32'h00068313;
mem['h158F] = 32'h00112623;
mem['h1590] = 32'h00060513;
mem['h1591] = 32'h000E0893;
mem['h1592] = 32'h00060693;
mem['h1593] = 32'h00000713;
mem['h1594] = 32'h00000793;
mem['h1595] = 32'h00000813;
mem['h1596] = 32'h0016FE93;
mem['h1597] = 32'h00171613;
mem['h1598] = 32'h000E8A63;
mem['h1599] = 32'h01088833;
mem['h159A] = 32'h00E787B3;
mem['h159B] = 32'h01183733;
mem['h159C] = 32'h00F707B3;
mem['h159D] = 32'h01F8D713;
mem['h159E] = 32'h0016D693;
mem['h159F] = 32'h00E66733;
mem['h15A0] = 32'h00189893;
mem['h15A1] = 32'hFC069AE3;
mem['h15A2] = 32'h00058663;
mem['h15A3] = 32'hF81FF0EF;
mem['h15A4] = 32'h00A787B3;
mem['h15A5] = 32'h00030A63;
mem['h15A6] = 32'h000E0513;
mem['h15A7] = 32'h00030593;
mem['h15A8] = 32'hF6DFF0EF;
mem['h15A9] = 32'h00F507B3;
mem['h15AA] = 32'h00C12083;
mem['h15AB] = 32'h00080513;
mem['h15AC] = 32'h00078593;
mem['h15AD] = 32'h01010113;
mem['h15AE] = 32'h00008067;
mem['h15AF] = 32'h06054063;
mem['h15B0] = 32'h0605C663;
mem['h15B1] = 32'h00058613;
mem['h15B2] = 32'h00050593;
mem['h15B3] = 32'hFFF00513;
mem['h15B4] = 32'h02060C63;
mem['h15B5] = 32'h00100693;
mem['h15B6] = 32'h00B67A63;
mem['h15B7] = 32'h00C05863;
mem['h15B8] = 32'h00161613;
mem['h15B9] = 32'h00169693;
mem['h15BA] = 32'hFEB66AE3;
mem['h15BB] = 32'h00000513;
mem['h15BC] = 32'h00C5E663;
mem['h15BD] = 32'h40C585B3;
mem['h15BE] = 32'h00D56533;
mem['h15BF] = 32'h0016D693;
mem['h15C0] = 32'h00165613;
mem['h15C1] = 32'hFE0696E3;
mem['h15C2] = 32'h00008067;
mem['h15C3] = 32'h00008293;
mem['h15C4] = 32'hFB5FF0EF;
mem['h15C5] = 32'h00058513;
mem['h15C6] = 32'h00028067;
mem['h15C7] = 32'h40A00533;
mem['h15C8] = 32'h00B04863;
mem['h15C9] = 32'h40B005B3;
mem['h15CA] = 32'hF9DFF06F;
mem['h15CB] = 32'h40B005B3;
mem['h15CC] = 32'h00008293;
mem['h15CD] = 32'hF91FF0EF;
mem['h15CE] = 32'h40A00533;
mem['h15CF] = 32'h00028067;
mem['h15D0] = 32'h00008293;
mem['h15D1] = 32'h0005CA63;
mem['h15D2] = 32'h00054C63;
mem['h15D3] = 32'hF79FF0EF;
mem['h15D4] = 32'h00058513;
mem['h15D5] = 32'h00028067;
mem['h15D6] = 32'h40B005B3;
mem['h15D7] = 32'hFE0558E3;
mem['h15D8] = 32'h40A00533;
mem['h15D9] = 32'hF61FF0EF;
mem['h15DA] = 32'h40B00533;
mem['h15DB] = 32'h00028067;
mem['h15DC] = 32'h33323130;
mem['h15DD] = 32'h37363534;
mem['h15DE] = 32'h42413938;
mem['h15DF] = 32'h46454443;
mem['h15E0] = 32'h00000000;
mem['h15E1] = 32'h00282020;
mem['h15E2] = 32'h50492029;
mem['h15E3] = 32'h0000203A;
mem['h15E4] = 32'h614D202C;
mem['h15E5] = 32'h203A6B73;
mem['h15E6] = 32'h00000000;
mem['h15E7] = 32'h6550202C;
mem['h15E8] = 32'h69207265;
mem['h15E9] = 32'h7865646E;
mem['h15EA] = 32'h0000203A;
mem['h15EB] = 32'h7344202C;
mem['h15EC] = 32'h00203A74;
mem['h15ED] = 32'h6F4C2029;
mem['h15EE] = 32'h206C6163;
mem['h15EF] = 32'h3A43414D;
mem['h15F0] = 32'h00000020;
mem['h15F1] = 32'h6F4C202C;
mem['h15F2] = 32'h206C6163;
mem['h15F3] = 32'h203A5049;
mem['h15F4] = 32'h00000000;
mem['h15F5] = 32'h6F4C202C;
mem['h15F6] = 32'h206C6163;
mem['h15F7] = 32'h74726F70;
mem['h15F8] = 32'h0000203A;
mem['h15F9] = 32'h6F4C202C;
mem['h15FA] = 32'h206C6163;
mem['h15FB] = 32'h203A4449;
mem['h15FC] = 32'h00007830;
mem['h15FD] = 32'h20200A0D;
mem['h15FE] = 32'h65522020;
mem['h15FF] = 32'h65746F6D;
mem['h1600] = 32'h43414D20;
mem['h1601] = 32'h0000203A;
mem['h1602] = 32'h6552202C;
mem['h1603] = 32'h65746F6D;
mem['h1604] = 32'h3A504920;
mem['h1605] = 32'h00000020;
mem['h1606] = 32'h6552202C;
mem['h1607] = 32'h65746F6D;
mem['h1608] = 32'h726F7020;
mem['h1609] = 32'h00203A74;
mem['h160A] = 32'h6552202C;
mem['h160B] = 32'h65746F6D;
mem['h160C] = 32'h3A444920;
mem['h160D] = 32'h00783020;
mem['h160E] = 32'h20200A0D;
mem['h160F] = 32'h6E452020;
mem['h1610] = 32'h70797263;
mem['h1611] = 32'h6E6F6974;
mem['h1612] = 32'h79656B20;
mem['h1613] = 32'h7830203A;
mem['h1614] = 32'h00000000;
mem['h1615] = 32'h20200A0D;
mem['h1616] = 32'h65442020;
mem['h1617] = 32'h70797263;
mem['h1618] = 32'h6E6F6974;
mem['h1619] = 32'h79656B20;
mem['h161A] = 32'h7830203A;
mem['h161B] = 32'h00000000;
mem['h161C] = 32'h20200A0D;
mem['h161D] = 32'h65532020;
mem['h161E] = 32'h6320646E;
mem['h161F] = 32'h746E756F;
mem['h1620] = 32'h203A7265;
mem['h1621] = 32'h00007830;
mem['h1622] = 32'h20200A0D;
mem['h1623] = 32'h65522020;
mem['h1624] = 32'h63207663;
mem['h1625] = 32'h746E756F;
mem['h1626] = 32'h203A7265;
mem['h1627] = 32'h00007830;
mem['h1628] = 32'h7774654E;
mem['h1629] = 32'h206B726F;
mem['h162A] = 32'h666E6F63;
mem['h162B] = 32'h72756769;
mem['h162C] = 32'h6F697461;
mem['h162D] = 32'h0A0D3A6E;
mem['h162E] = 32'h00000000;
mem['h162F] = 32'h50492020;
mem['h1630] = 32'h64646120;
mem['h1631] = 32'h73736572;
mem['h1632] = 32'h2020203A;
mem['h1633] = 32'h20202020;
mem['h1634] = 32'h00000020;
mem['h1635] = 32'h20200A0D;
mem['h1636] = 32'h6E627553;
mem['h1637] = 32'h6D207465;
mem['h1638] = 32'h3A6B7361;
mem['h1639] = 32'h20202020;
mem['h163A] = 32'h00202020;
mem['h163B] = 32'h20200A0D;
mem['h163C] = 32'h2043414D;
mem['h163D] = 32'h72646461;
mem['h163E] = 32'h3A737365;
mem['h163F] = 32'h20202020;
mem['h1640] = 32'h00202020;
mem['h1641] = 32'h20200A0D;
mem['h1642] = 32'h61666544;
mem['h1643] = 32'h20746C75;
mem['h1644] = 32'h65746167;
mem['h1645] = 32'h3A796177;
mem['h1646] = 32'h00202020;
mem['h1647] = 32'h20200A0D;
mem['h1648] = 32'h61666544;
mem['h1649] = 32'h20746C75;
mem['h164A] = 32'h65746E69;
mem['h164B] = 32'h63616672;
mem['h164C] = 32'h00203A65;
mem['h164D] = 32'h69646441;
mem['h164E] = 32'h6E6F6974;
mem['h164F] = 32'h61206C61;
mem['h1650] = 32'h65687475;
mem['h1651] = 32'h6369746E;
mem['h1652] = 32'h64657461;
mem['h1653] = 32'h74616420;
mem['h1654] = 32'h00000061;
mem['h1655] = 32'h6C6C6548;
mem['h1656] = 32'h4843206F;
mem['h1657] = 32'h43494C49;
mem['h1658] = 32'h73706968;
mem['h1659] = 32'h57202D20;
mem['h165A] = 32'h67657269;
mem['h165B] = 32'h64726175;
mem['h165C] = 32'h61657420;
mem['h165D] = 32'h6C202C6D;
mem['h165E] = 32'h73277465;
mem['h165F] = 32'h73657420;
mem['h1660] = 32'h68742074;
mem['h1661] = 32'h61207369;
mem['h1662] = 32'h21646165;
mem['h1663] = 32'h00000000;
mem['h1664] = 32'h43616843;
mem['h1665] = 32'h30326168;
mem['h1666] = 32'h6C6F502D;
mem['h1667] = 32'h30333179;
mem['h1668] = 32'h65742035;
mem['h1669] = 32'h70207473;
mem['h166A] = 32'h65737361;
mem['h166B] = 32'h0A0D2164;
mem['h166C] = 32'h00000000;
mem['h166D] = 32'h43616843;
mem['h166E] = 32'h30326168;
mem['h166F] = 32'h6C6F502D;
mem['h1670] = 32'h30333179;
mem['h1671] = 32'h65742035;
mem['h1672] = 32'h66207473;
mem['h1673] = 32'h656C6961;
mem['h1674] = 32'h0A0D2164;
mem['h1675] = 32'h00000000;
mem['h1676] = 32'h83828180;
mem['h1677] = 32'h87868584;
mem['h1678] = 32'h8B8A8988;
mem['h1679] = 32'h8F8E8D8C;
mem['h167A] = 32'h93929190;
mem['h167B] = 32'h97969594;
mem['h167C] = 32'h9B9A9998;
mem['h167D] = 32'h9F9E9D9C;
mem['h167E] = 32'h00000000;
mem['h167F] = 32'h61480A0D;
mem['h1680] = 32'h61776472;
mem['h1681] = 32'h49206572;
mem['h1682] = 32'h696D2044;
mem['h1683] = 32'h74616D73;
mem['h1684] = 32'h20216863;
mem['h1685] = 32'h746C6148;
mem['h1686] = 32'h2E676E69;
mem['h1687] = 32'h0A0D2E2E;
mem['h1688] = 32'h00000000;
mem['h1689] = 32'h3D3D0A0D;
mem['h168A] = 32'h3D3D3D3D;
mem['h168B] = 32'h3D3D3D3D;
mem['h168C] = 32'h3D3D3D3D;
mem['h168D] = 32'h3D3D3D3D;
mem['h168E] = 32'h3D3D3D3D;
mem['h168F] = 32'h3D3D3D3D;
mem['h1690] = 32'h3D3D3D3D;
mem['h1691] = 32'h3D3D3D3D;
mem['h1692] = 32'h3D3D3D3D;
mem['h1693] = 32'h3D3D3D3D;
mem['h1694] = 32'h00000A0D;
mem['h1695] = 32'h20202020;
mem['h1696] = 32'h20202020;
mem['h1697] = 32'h69572020;
mem['h1698] = 32'h75476572;
mem['h1699] = 32'h20647261;
mem['h169A] = 32'h41475046;
mem['h169B] = 32'h00007620;
mem['h169C] = 32'h20200A0D;
mem['h169D] = 32'h706F4320;
mem['h169E] = 32'h67697279;
mem['h169F] = 32'hC2207468;
mem['h16A0] = 32'h303220A9;
mem['h16A1] = 32'h322D3432;
mem['h16A2] = 32'h20363230;
mem['h16A3] = 32'h6C696843;
mem['h16A4] = 32'h48432E69;
mem['h16A5] = 32'h2A535049;
mem['h16A6] = 32'h0A0D6162;
mem['h16A7] = 32'h00000000;
mem['h16A8] = 32'h3D3D3D3D;
mem['h16A9] = 32'h3D3D3D3D;
mem['h16AA] = 32'h3D3D3D3D;
mem['h16AB] = 32'h3D3D3D3D;
mem['h16AC] = 32'h3D3D3D3D;
mem['h16AD] = 32'h3D3D3D3D;
mem['h16AE] = 32'h3D3D3D3D;
mem['h16AF] = 32'h3D3D3D3D;
mem['h16B0] = 32'h3D3D3D3D;
mem['h16B1] = 32'h3D3D3D3D;
mem['h16B2] = 32'h0A0D3D3D;
mem['h16B3] = 32'h00000000;
mem['h16B4] = 32'h746F6F42;
mem['h16B5] = 32'h20676E69;
mem['h16B6] = 32'h2E2E7075;
mem['h16B7] = 32'h000A0D2E;
mem['h16B8] = 32'h79540A0D;
mem['h16B9] = 32'h27206570;
mem['h16BA] = 32'h706C6568;
mem['h16BB] = 32'h6F742027;
mem['h16BC] = 32'h73696420;
mem['h16BD] = 32'h79616C70;
mem['h16BE] = 32'h6D6F6320;
mem['h16BF] = 32'h646E616D;
mem['h16C0] = 32'h0A0D2E73;
mem['h16C1] = 32'h00000000;
mem['h16C2] = 32'h72697728;
mem['h16C3] = 32'h61756765;
mem['h16C4] = 32'h662D6472;
mem['h16C5] = 32'h29616770;
mem['h16C6] = 32'h00002023;
mem['h16C7] = 32'h4E203C3C;
mem['h16C8] = 32'h505F5445;
mem['h16C9] = 32'h4F544F52;
mem['h16CA] = 32'h4B4E555F;
mem['h16CB] = 32'h4E574F4E;
mem['h16CC] = 32'h0000203A;
mem['h16CD] = 32'h4E203C3C;
mem['h16CE] = 32'h505F5445;
mem['h16CF] = 32'h4F544F52;
mem['h16D0] = 32'h5052415F;
mem['h16D1] = 32'h0000203A;
mem['h16D2] = 32'h4E203E3E;
mem['h16D3] = 32'h505F5445;
mem['h16D4] = 32'h4F544F52;
mem['h16D5] = 32'h5052415F;
mem['h16D6] = 32'h0000203A;
mem['h16D7] = 32'h4E203C3C;
mem['h16D8] = 32'h505F5445;
mem['h16D9] = 32'h4F544F52;
mem['h16DA] = 32'h4D43495F;
mem['h16DB] = 32'h00203A50;
mem['h16DC] = 32'h4E203E3E;
mem['h16DD] = 32'h505F5445;
mem['h16DE] = 32'h4F544F52;
mem['h16DF] = 32'h4D43495F;
mem['h16E0] = 32'h00203A50;
mem['h16E1] = 32'h4E203C3C;
mem['h16E2] = 32'h505F5445;
mem['h16E3] = 32'h4F544F52;
mem['h16E4] = 32'h5044555F;
mem['h16E5] = 32'h0000203A;
mem['h16E6] = 32'h74736574;
mem['h16E7] = 32'h61686320;
mem['h16E8] = 32'h32616863;
mem['h16E9] = 32'h6C6F7030;
mem['h16EA] = 32'h30333179;
mem['h16EB] = 32'h00000A35;
mem['h16EC] = 32'h74736574;
mem['h16ED] = 32'h616C6220;
mem['h16EE] = 32'h7332656B;
mem['h16EF] = 32'h0000000A;
mem['h16F0] = 32'h00636261;
mem['h16F1] = 32'h4B414C42;
mem['h16F2] = 32'h20733245;
mem['h16F3] = 32'h74736574;
mem['h16F4] = 32'h73617020;
mem['h16F5] = 32'h21646573;
mem['h16F6] = 32'h00000A0D;
mem['h16F7] = 32'h4B414C42;
mem['h16F8] = 32'h20733245;
mem['h16F9] = 32'h74736574;
mem['h16FA] = 32'h69616620;
mem['h16FB] = 32'h2164656C;
mem['h16FC] = 32'h00000A0D;
mem['h16FD] = 32'h74736574;
mem['h16FE] = 32'h72756320;
mem['h16FF] = 32'h35326576;
mem['h1700] = 32'h0A393135;
mem['h1701] = 32'h00000000;
mem['h1702] = 32'h2079654B;
mem['h1703] = 32'h68637865;
mem['h1704] = 32'h65676E61;
mem['h1705] = 32'h63757320;
mem['h1706] = 32'h73736563;
mem['h1707] = 32'h216C7566;
mem['h1708] = 32'h696C4120;
mem['h1709] = 32'h61206563;
mem['h170A] = 32'h4220646E;
mem['h170B] = 32'h6820626F;
mem['h170C] = 32'h20657661;
mem['h170D] = 32'h20656874;
mem['h170E] = 32'h656D6173;
mem['h170F] = 32'h61687320;
mem['h1710] = 32'h20646572;
mem['h1711] = 32'h72636573;
mem['h1712] = 32'h0A0D7465;
mem['h1713] = 32'h00000000;
mem['h1714] = 32'h2079654B;
mem['h1715] = 32'h68637865;
mem['h1716] = 32'h65676E61;
mem['h1717] = 32'h69616620;
mem['h1718] = 32'h2164656C;
mem['h1719] = 32'h61685320;
mem['h171A] = 32'h20646572;
mem['h171B] = 32'h72636573;
mem['h171C] = 32'h20737465;
mem['h171D] = 32'h276E6F64;
mem['h171E] = 32'h616D2074;
mem['h171F] = 32'h2E686374;
mem['h1720] = 32'h00000A0D;
mem['h1721] = 32'h74736574;
mem['h1722] = 32'h676E7220;
mem['h1723] = 32'h0000000A;
mem['h1724] = 32'h656E6547;
mem['h1725] = 32'h69746172;
mem['h1726] = 32'h7220676E;
mem['h1727] = 32'h6F646E61;
mem['h1728] = 32'h3233206D;
mem['h1729] = 32'h74796220;
mem['h172A] = 32'h203A7365;
mem['h172B] = 32'h00000000;
mem['h172C] = 32'h656E6547;
mem['h172D] = 32'h69746172;
mem['h172E] = 32'h7220676E;
mem['h172F] = 32'h6F646E61;
mem['h1730] = 32'h756E206D;
mem['h1731] = 32'h7265626D;
mem['h1732] = 32'h74656220;
mem['h1733] = 32'h6E656577;
mem['h1734] = 32'h20303120;
mem['h1735] = 32'h20646E61;
mem['h1736] = 32'h30303031;
mem['h1737] = 32'h0000203A;
mem['h1738] = 32'h74736574;
mem['h1739] = 32'h6D697420;
mem['h173A] = 32'h000A7265;
mem['h173B] = 32'h0000002E;
mem['h173C] = 32'h65540A0D;
mem['h173D] = 32'h70207473;
mem['h173E] = 32'h65737361;
mem['h173F] = 32'h0A0D2164;
mem['h1740] = 32'h00000000;
mem['h1741] = 32'h776F6873;
mem['h1742] = 32'h74656E20;
mem['h1743] = 32'h6B726F77;
mem['h1744] = 32'h0000000A;
mem['h1745] = 32'h666E6F63;
mem['h1746] = 32'h6E206769;
mem['h1747] = 32'h6F777465;
mem['h1748] = 32'h000A6B72;
mem['h1749] = 32'h65746E45;
mem['h174A] = 32'h656E2072;
mem['h174B] = 32'h656E2077;
mem['h174C] = 32'h726F7774;
mem['h174D] = 32'h6F63206B;
mem['h174E] = 32'h6769666E;
mem['h174F] = 32'h74617275;
mem['h1750] = 32'h3A6E6F69;
mem['h1751] = 32'h00000A0D;
mem['h1752] = 32'h50492020;
mem['h1753] = 32'h64646120;
mem['h1754] = 32'h73736572;
mem['h1755] = 32'h00005B20;
mem['h1756] = 32'h75532020;
mem['h1757] = 32'h74656E62;
mem['h1758] = 32'h73616D20;
mem['h1759] = 32'h005B206B;
mem['h175A] = 32'h65472020;
mem['h175B] = 32'h6172656E;
mem['h175C] = 32'h6E206574;
mem['h175D] = 32'h4D207765;
mem['h175E] = 32'h61204341;
mem['h175F] = 32'h65726464;
mem['h1760] = 32'h203F7373;
mem['h1761] = 32'h6E2F7928;
mem['h1762] = 32'h6E5B2029;
mem['h1763] = 32'h00203A5D;
mem['h1764] = 32'h65442020;
mem['h1765] = 32'h6C756166;
mem['h1766] = 32'h61672074;
mem['h1767] = 32'h61776574;
mem['h1768] = 32'h005B2079;
mem['h1769] = 32'h65442020;
mem['h176A] = 32'h6C756166;
mem['h176B] = 32'h6E692074;
mem['h176C] = 32'h66726574;
mem['h176D] = 32'h20656361;
mem['h176E] = 32'h332D3028;
mem['h176F] = 32'h005B2029;
mem['h1770] = 32'h7774654E;
mem['h1771] = 32'h206B726F;
mem['h1772] = 32'h666E6F63;
mem['h1773] = 32'h72756769;
mem['h1774] = 32'h6F697461;
mem['h1775] = 32'h7075206E;
mem['h1776] = 32'h65746164;
mem['h1777] = 32'h0A0D2E64;
mem['h1778] = 32'h00000000;
mem['h1779] = 32'h776F6873;
mem['h177A] = 32'h756F7220;
mem['h177B] = 32'h0A736574;
mem['h177C] = 32'h00000000;
mem['h177D] = 32'h74756F52;
mem['h177E] = 32'h20676E69;
mem['h177F] = 32'h6C626174;
mem['h1780] = 32'h0A0D3A65;
mem['h1781] = 32'h00000000;
mem['h1782] = 32'h666E6F63;
mem['h1783] = 32'h72206769;
mem['h1784] = 32'h6574756F;
mem['h1785] = 32'h00000A73;
mem['h1786] = 32'h65746E45;
mem['h1787] = 32'h656E2072;
mem['h1788] = 32'h6F722077;
mem['h1789] = 32'h6E697475;
mem['h178A] = 32'h61742067;
mem['h178B] = 32'h20656C62;
mem['h178C] = 32'h72746E65;
mem['h178D] = 32'h0A0D3A79;
mem['h178E] = 32'h00000000;
mem['h178F] = 32'h6E452020;
mem['h1790] = 32'h20797274;
mem['h1791] = 32'h65646E69;
mem['h1792] = 32'h30282078;
mem['h1793] = 32'h2933362D;
mem['h1794] = 32'h5D305B20;
mem['h1795] = 32'h0000203A;
mem['h1796] = 32'h65442020;
mem['h1797] = 32'h6E697473;
mem['h1798] = 32'h6F697461;
mem['h1799] = 32'h5049206E;
mem['h179A] = 32'h64646120;
mem['h179B] = 32'h73736572;
mem['h179C] = 32'h00005B20;
mem['h179D] = 32'h65502020;
mem['h179E] = 32'h69207265;
mem['h179F] = 32'h7865646E;
mem['h17A0] = 32'h2D302820;
mem['h17A1] = 32'h20293336;
mem['h17A2] = 32'h0000005B;
mem['h17A3] = 32'h73442020;
mem['h17A4] = 32'h30282074;
mem['h17A5] = 32'h2029332D;
mem['h17A6] = 32'h0000005B;
mem['h17A7] = 32'h74756F52;
mem['h17A8] = 32'h20676E69;
mem['h17A9] = 32'h6C626174;
mem['h17AA] = 32'h6E652065;
mem['h17AB] = 32'h20797274;
mem['h17AC] = 32'h61647075;
mem['h17AD] = 32'h2E646574;
mem['h17AE] = 32'h00000A0D;
mem['h17AF] = 32'h776F6873;
mem['h17B0] = 32'h79726320;
mem['h17B1] = 32'h6B6F7470;
mem['h17B2] = 32'h0A737965;
mem['h17B3] = 32'h00000000;
mem['h17B4] = 32'h70797243;
mem['h17B5] = 32'h656B6F74;
mem['h17B6] = 32'h61742079;
mem['h17B7] = 32'h3A656C62;
mem['h17B8] = 32'h00000A0D;
mem['h17B9] = 32'h666E6F63;
mem['h17BA] = 32'h63206769;
mem['h17BB] = 32'h74707972;
mem['h17BC] = 32'h79656B6F;
mem['h17BD] = 32'h00000A73;
mem['h17BE] = 32'h65746E45;
mem['h17BF] = 32'h656E2072;
mem['h17C0] = 32'h72632077;
mem['h17C1] = 32'h6F747079;
mem['h17C2] = 32'h2079656B;
mem['h17C3] = 32'h6C626174;
mem['h17C4] = 32'h6E652065;
mem['h17C5] = 32'h3A797274;
mem['h17C6] = 32'h00000A0D;
mem['h17C7] = 32'h6F4C2020;
mem['h17C8] = 32'h206C6163;
mem['h17C9] = 32'h2043414D;
mem['h17CA] = 32'h72646461;
mem['h17CB] = 32'h20737365;
mem['h17CC] = 32'h0000005B;
mem['h17CD] = 32'h6F4C2020;
mem['h17CE] = 32'h206C6163;
mem['h17CF] = 32'h61205049;
mem['h17D0] = 32'h65726464;
mem['h17D1] = 32'h5B207373;
mem['h17D2] = 32'h00000000;
mem['h17D3] = 32'h6F4C2020;
mem['h17D4] = 32'h206C6163;
mem['h17D5] = 32'h74726F70;
mem['h17D6] = 32'h2D302820;
mem['h17D7] = 32'h33353536;
mem['h17D8] = 32'h5B202935;
mem['h17D9] = 32'h00000000;
mem['h17DA] = 32'h6F4C2020;
mem['h17DB] = 32'h206C6163;
mem['h17DC] = 32'h28204449;
mem['h17DD] = 32'h65682038;
mem['h17DE] = 32'h69642078;
mem['h17DF] = 32'h73746967;
mem['h17E0] = 32'h005B2029;
mem['h17E1] = 32'h65522020;
mem['h17E2] = 32'h65746F6D;
mem['h17E3] = 32'h43414D20;
mem['h17E4] = 32'h64646120;
mem['h17E5] = 32'h73736572;
mem['h17E6] = 32'h00005B20;
mem['h17E7] = 32'h65522020;
mem['h17E8] = 32'h65746F6D;
mem['h17E9] = 32'h20504920;
mem['h17EA] = 32'h72646461;
mem['h17EB] = 32'h20737365;
mem['h17EC] = 32'h0000005B;
mem['h17ED] = 32'h65522020;
mem['h17EE] = 32'h65746F6D;
mem['h17EF] = 32'h726F7020;
mem['h17F0] = 32'h30282074;
mem['h17F1] = 32'h3535362D;
mem['h17F2] = 32'h20293533;
mem['h17F3] = 32'h0000005B;
mem['h17F4] = 32'h65522020;
mem['h17F5] = 32'h65746F6D;
mem['h17F6] = 32'h20444920;
mem['h17F7] = 32'h68203828;
mem['h17F8] = 32'h64207865;
mem['h17F9] = 32'h74696769;
mem['h17FA] = 32'h5B202973;
mem['h17FB] = 32'h00000000;
mem['h17FC] = 32'h6E452020;
mem['h17FD] = 32'h70797263;
mem['h17FE] = 32'h6E6F6974;
mem['h17FF] = 32'h79656B20;
mem['h1800] = 32'h73312820;
mem['h1801] = 32'h20382074;
mem['h1802] = 32'h20786568;
mem['h1803] = 32'h69676964;
mem['h1804] = 32'h20297374;
mem['h1805] = 32'h0000005B;
mem['h1806] = 32'h6E452020;
mem['h1807] = 32'h70797263;
mem['h1808] = 32'h6E6F6974;
mem['h1809] = 32'h79656B20;
mem['h180A] = 32'h6E322820;
mem['h180B] = 32'h20382064;
mem['h180C] = 32'h20786568;
mem['h180D] = 32'h69676964;
mem['h180E] = 32'h20297374;
mem['h180F] = 32'h0000005B;
mem['h1810] = 32'h6E452020;
mem['h1811] = 32'h70797263;
mem['h1812] = 32'h6E6F6974;
mem['h1813] = 32'h79656B20;
mem['h1814] = 32'h72332820;
mem['h1815] = 32'h20382064;
mem['h1816] = 32'h20786568;
mem['h1817] = 32'h69676964;
mem['h1818] = 32'h20297374;
mem['h1819] = 32'h0000005B;
mem['h181A] = 32'h6E452020;
mem['h181B] = 32'h70797263;
mem['h181C] = 32'h6E6F6974;
mem['h181D] = 32'h79656B20;
mem['h181E] = 32'h74342820;
mem['h181F] = 32'h20382068;
mem['h1820] = 32'h20786568;
mem['h1821] = 32'h69676964;
mem['h1822] = 32'h20297374;
mem['h1823] = 32'h0000005B;
mem['h1824] = 32'h6E452020;
mem['h1825] = 32'h70797263;
mem['h1826] = 32'h6E6F6974;
mem['h1827] = 32'h79656B20;
mem['h1828] = 32'h74352820;
mem['h1829] = 32'h20382068;
mem['h182A] = 32'h20786568;
mem['h182B] = 32'h69676964;
mem['h182C] = 32'h20297374;
mem['h182D] = 32'h0000005B;
mem['h182E] = 32'h6E452020;
mem['h182F] = 32'h70797263;
mem['h1830] = 32'h6E6F6974;
mem['h1831] = 32'h79656B20;
mem['h1832] = 32'h74362820;
mem['h1833] = 32'h20382068;
mem['h1834] = 32'h20786568;
mem['h1835] = 32'h69676964;
mem['h1836] = 32'h20297374;
mem['h1837] = 32'h0000005B;
mem['h1838] = 32'h6E452020;
mem['h1839] = 32'h70797263;
mem['h183A] = 32'h6E6F6974;
mem['h183B] = 32'h79656B20;
mem['h183C] = 32'h74372820;
mem['h183D] = 32'h20382068;
mem['h183E] = 32'h20786568;
mem['h183F] = 32'h69676964;
mem['h1840] = 32'h20297374;
mem['h1841] = 32'h0000005B;
mem['h1842] = 32'h6E452020;
mem['h1843] = 32'h70797263;
mem['h1844] = 32'h6E6F6974;
mem['h1845] = 32'h79656B20;
mem['h1846] = 32'h74382820;
mem['h1847] = 32'h20382068;
mem['h1848] = 32'h20786568;
mem['h1849] = 32'h69676964;
mem['h184A] = 32'h20297374;
mem['h184B] = 32'h0000005B;
mem['h184C] = 32'h65442020;
mem['h184D] = 32'h70797263;
mem['h184E] = 32'h6E6F6974;
mem['h184F] = 32'h79656B20;
mem['h1850] = 32'h73312820;
mem['h1851] = 32'h20382074;
mem['h1852] = 32'h20786568;
mem['h1853] = 32'h69676964;
mem['h1854] = 32'h20297374;
mem['h1855] = 32'h0000005B;
mem['h1856] = 32'h65442020;
mem['h1857] = 32'h70797263;
mem['h1858] = 32'h6E6F6974;
mem['h1859] = 32'h79656B20;
mem['h185A] = 32'h6E322820;
mem['h185B] = 32'h20382064;
mem['h185C] = 32'h20786568;
mem['h185D] = 32'h69676964;
mem['h185E] = 32'h20297374;
mem['h185F] = 32'h0000005B;
mem['h1860] = 32'h65442020;
mem['h1861] = 32'h70797263;
mem['h1862] = 32'h6E6F6974;
mem['h1863] = 32'h79656B20;
mem['h1864] = 32'h72332820;
mem['h1865] = 32'h20382064;
mem['h1866] = 32'h20786568;
mem['h1867] = 32'h69676964;
mem['h1868] = 32'h20297374;
mem['h1869] = 32'h0000005B;
mem['h186A] = 32'h65442020;
mem['h186B] = 32'h70797263;
mem['h186C] = 32'h6E6F6974;
mem['h186D] = 32'h79656B20;
mem['h186E] = 32'h74342820;
mem['h186F] = 32'h20382068;
mem['h1870] = 32'h20786568;
mem['h1871] = 32'h69676964;
mem['h1872] = 32'h20297374;
mem['h1873] = 32'h0000005B;
mem['h1874] = 32'h65442020;
mem['h1875] = 32'h70797263;
mem['h1876] = 32'h6E6F6974;
mem['h1877] = 32'h79656B20;
mem['h1878] = 32'h74352820;
mem['h1879] = 32'h20382068;
mem['h187A] = 32'h20786568;
mem['h187B] = 32'h69676964;
mem['h187C] = 32'h20297374;
mem['h187D] = 32'h0000005B;
mem['h187E] = 32'h65442020;
mem['h187F] = 32'h70797263;
mem['h1880] = 32'h6E6F6974;
mem['h1881] = 32'h79656B20;
mem['h1882] = 32'h74362820;
mem['h1883] = 32'h20382068;
mem['h1884] = 32'h20786568;
mem['h1885] = 32'h69676964;
mem['h1886] = 32'h20297374;
mem['h1887] = 32'h0000005B;
mem['h1888] = 32'h65442020;
mem['h1889] = 32'h70797263;
mem['h188A] = 32'h6E6F6974;
mem['h188B] = 32'h79656B20;
mem['h188C] = 32'h74372820;
mem['h188D] = 32'h20382068;
mem['h188E] = 32'h20786568;
mem['h188F] = 32'h69676964;
mem['h1890] = 32'h20297374;
mem['h1891] = 32'h0000005B;
mem['h1892] = 32'h65442020;
mem['h1893] = 32'h70797263;
mem['h1894] = 32'h6E6F6974;
mem['h1895] = 32'h79656B20;
mem['h1896] = 32'h74382820;
mem['h1897] = 32'h20382068;
mem['h1898] = 32'h20786568;
mem['h1899] = 32'h69676964;
mem['h189A] = 32'h20297374;
mem['h189B] = 32'h0000005B;
mem['h189C] = 32'h65522020;
mem['h189D] = 32'h20746573;
mem['h189E] = 32'h646E6573;
mem['h189F] = 32'h6365722F;
mem['h18A0] = 32'h6F632076;
mem['h18A1] = 32'h65746E75;
mem['h18A2] = 32'h203F7372;
mem['h18A3] = 32'h6E2F7928;
mem['h18A4] = 32'h6E5B2029;
mem['h18A5] = 32'h00203A5D;
mem['h18A6] = 32'h70797243;
mem['h18A7] = 32'h656B6F74;
mem['h18A8] = 32'h61742079;
mem['h18A9] = 32'h20656C62;
mem['h18AA] = 32'h72746E65;
mem['h18AB] = 32'h70752079;
mem['h18AC] = 32'h65746164;
mem['h18AD] = 32'h0A0D2E64;
mem['h18AE] = 32'h00000000;
mem['h18AF] = 32'h75626564;
mem['h18B0] = 32'h00000A67;
mem['h18B1] = 32'h75626544;
mem['h18B2] = 32'h6F6D2067;
mem['h18B3] = 32'h00206564;
mem['h18B4] = 32'h62616E65;
mem['h18B5] = 32'h2E64656C;
mem['h18B6] = 32'h00000A0D;
mem['h18B7] = 32'h61736964;
mem['h18B8] = 32'h64656C62;
mem['h18B9] = 32'h000A0D2E;
mem['h18BA] = 32'h6F626572;
mem['h18BB] = 32'h000A746F;
mem['h18BC] = 32'h706C6568;
mem['h18BD] = 32'h0000000A;
mem['h18BE] = 32'h69617641;
mem['h18BF] = 32'h6C62616C;
mem['h18C0] = 32'h6F632065;
mem['h18C1] = 32'h6E616D6D;
mem['h18C2] = 32'h0D3A7364;
mem['h18C3] = 32'h0000000A;
mem['h18C4] = 32'h65742020;
mem['h18C5] = 32'h63207473;
mem['h18C6] = 32'h68636168;
mem['h18C7] = 32'h70303261;
mem['h18C8] = 32'h31796C6F;
mem['h18C9] = 32'h20353033;
mem['h18CA] = 32'h54202D20;
mem['h18CB] = 32'h20747365;
mem['h18CC] = 32'h43616843;
mem['h18CD] = 32'h30326168;
mem['h18CE] = 32'h6C6F502D;
mem['h18CF] = 32'h30333179;
mem['h18D0] = 32'h45412035;
mem['h18D1] = 32'h0A0D4441;
mem['h18D2] = 32'h00000000;
mem['h18D3] = 32'h65742020;
mem['h18D4] = 32'h62207473;
mem['h18D5] = 32'h656B616C;
mem['h18D6] = 32'h20207332;
mem['h18D7] = 32'h20202020;
mem['h18D8] = 32'h20202020;
mem['h18D9] = 32'h54202D20;
mem['h18DA] = 32'h20747365;
mem['h18DB] = 32'h4B414C42;
mem['h18DC] = 32'h20733245;
mem['h18DD] = 32'h68736168;
mem['h18DE] = 32'h6E756620;
mem['h18DF] = 32'h6F697463;
mem['h18E0] = 32'h000A0D6E;
mem['h18E1] = 32'h65742020;
mem['h18E2] = 32'h63207473;
mem['h18E3] = 32'h65767275;
mem['h18E4] = 32'h31353532;
mem['h18E5] = 32'h20202039;
mem['h18E6] = 32'h20202020;
mem['h18E7] = 32'h54202D20;
mem['h18E8] = 32'h20747365;
mem['h18E9] = 32'h76727543;
mem['h18EA] = 32'h35353265;
mem['h18EB] = 32'h6B203931;
mem['h18EC] = 32'h65207965;
mem['h18ED] = 32'h61686378;
mem['h18EE] = 32'h0D65676E;
mem['h18EF] = 32'h0000000A;
mem['h18F0] = 32'h65742020;
mem['h18F1] = 32'h72207473;
mem['h18F2] = 32'h2020676E;
mem['h18F3] = 32'h20202020;
mem['h18F4] = 32'h20202020;
mem['h18F5] = 32'h20202020;
mem['h18F6] = 32'h54202D20;
mem['h18F7] = 32'h20747365;
mem['h18F8] = 32'h646E6172;
mem['h18F9] = 32'h6E206D6F;
mem['h18FA] = 32'h65626D75;
mem['h18FB] = 32'h65672072;
mem['h18FC] = 32'h6172656E;
mem['h18FD] = 32'h0D726F74;
mem['h18FE] = 32'h0000000A;
mem['h18FF] = 32'h65742020;
mem['h1900] = 32'h74207473;
mem['h1901] = 32'h72656D69;
mem['h1902] = 32'h20202020;
mem['h1903] = 32'h20202020;
mem['h1904] = 32'h20202020;
mem['h1905] = 32'h54202D20;
mem['h1906] = 32'h20747365;
mem['h1907] = 32'h656D6974;
mem['h1908] = 32'h75662072;
mem['h1909] = 32'h6974636E;
mem['h190A] = 32'h6C616E6F;
mem['h190B] = 32'h0D797469;
mem['h190C] = 32'h0000000A;
mem['h190D] = 32'h68732020;
mem['h190E] = 32'h6E20776F;
mem['h190F] = 32'h6F777465;
mem['h1910] = 32'h20206B72;
mem['h1911] = 32'h20202020;
mem['h1912] = 32'h20202020;
mem['h1913] = 32'h53202D20;
mem['h1914] = 32'h20776F68;
mem['h1915] = 32'h7774656E;
mem['h1916] = 32'h206B726F;
mem['h1917] = 32'h666E6F63;
mem['h1918] = 32'h72756769;
mem['h1919] = 32'h6F697461;
mem['h191A] = 32'h000A0D6E;
mem['h191B] = 32'h6F632020;
mem['h191C] = 32'h6769666E;
mem['h191D] = 32'h74656E20;
mem['h191E] = 32'h6B726F77;
mem['h191F] = 32'h20202020;
mem['h1920] = 32'h20202020;
mem['h1921] = 32'h43202D20;
mem['h1922] = 32'h69666E6F;
mem['h1923] = 32'h65727567;
mem['h1924] = 32'h74656E20;
mem['h1925] = 32'h6B726F77;
mem['h1926] = 32'h74657320;
mem['h1927] = 32'h676E6974;
mem['h1928] = 32'h000A0D73;
mem['h1929] = 32'h68732020;
mem['h192A] = 32'h7220776F;
mem['h192B] = 32'h6574756F;
mem['h192C] = 32'h20202073;
mem['h192D] = 32'h20202020;
mem['h192E] = 32'h20202020;
mem['h192F] = 32'h53202D20;
mem['h1930] = 32'h20776F68;
mem['h1931] = 32'h74756F72;
mem['h1932] = 32'h20676E69;
mem['h1933] = 32'h6C626174;
mem['h1934] = 32'h000A0D65;
mem['h1935] = 32'h6F632020;
mem['h1936] = 32'h6769666E;
mem['h1937] = 32'h756F7220;
mem['h1938] = 32'h20736574;
mem['h1939] = 32'h20202020;
mem['h193A] = 32'h20202020;
mem['h193B] = 32'h43202D20;
mem['h193C] = 32'h69666E6F;
mem['h193D] = 32'h65727567;
mem['h193E] = 32'h756F7220;
mem['h193F] = 32'h676E6974;
mem['h1940] = 32'h62617420;
mem['h1941] = 32'h6520656C;
mem['h1942] = 32'h7972746E;
mem['h1943] = 32'h00000A0D;
mem['h1944] = 32'h68732020;
mem['h1945] = 32'h6320776F;
mem['h1946] = 32'h74707972;
mem['h1947] = 32'h79656B6F;
mem['h1948] = 32'h20202073;
mem['h1949] = 32'h20202020;
mem['h194A] = 32'h53202D20;
mem['h194B] = 32'h20776F68;
mem['h194C] = 32'h70797263;
mem['h194D] = 32'h656B6F74;
mem['h194E] = 32'h61742079;
mem['h194F] = 32'h0D656C62;
mem['h1950] = 32'h0000000A;
mem['h1951] = 32'h6F632020;
mem['h1952] = 32'h6769666E;
mem['h1953] = 32'h79726320;
mem['h1954] = 32'h6B6F7470;
mem['h1955] = 32'h20737965;
mem['h1956] = 32'h20202020;
mem['h1957] = 32'h43202D20;
mem['h1958] = 32'h69666E6F;
mem['h1959] = 32'h65727567;
mem['h195A] = 32'h79726320;
mem['h195B] = 32'h6B6F7470;
mem['h195C] = 32'h74207965;
mem['h195D] = 32'h656C6261;
mem['h195E] = 32'h746E6520;
mem['h195F] = 32'h0A0D7972;
mem['h1960] = 32'h00000000;
mem['h1961] = 32'h65642020;
mem['h1962] = 32'h20677562;
mem['h1963] = 32'h20202020;
mem['h1964] = 32'h20202020;
mem['h1965] = 32'h20202020;
mem['h1966] = 32'h20202020;
mem['h1967] = 32'h54202D20;
mem['h1968] = 32'h6C67676F;
mem['h1969] = 32'h65642065;
mem['h196A] = 32'h20677562;
mem['h196B] = 32'h65646F6D;
mem['h196C] = 32'h00000A0D;
mem['h196D] = 32'h65722020;
mem['h196E] = 32'h746F6F62;
mem['h196F] = 32'h20202020;
mem['h1970] = 32'h20202020;
mem['h1971] = 32'h20202020;
mem['h1972] = 32'h20202020;
mem['h1973] = 32'h52202D20;
mem['h1974] = 32'h6F6F6265;
mem['h1975] = 32'h68742074;
mem['h1976] = 32'h79732065;
mem['h1977] = 32'h6D657473;
mem['h1978] = 32'h00000A0D;
mem['h1979] = 32'h65682020;
mem['h197A] = 32'h2020706C;
mem['h197B] = 32'h20202020;
mem['h197C] = 32'h20202020;
mem['h197D] = 32'h20202020;
mem['h197E] = 32'h20202020;
mem['h197F] = 32'h53202D20;
mem['h1980] = 32'h20776F68;
mem['h1981] = 32'h73696874;
mem['h1982] = 32'h6C656820;
mem['h1983] = 32'h656D2070;
mem['h1984] = 32'h67617373;
mem['h1985] = 32'h000A0D65;
mem['h1986] = 32'h6E6B6E55;
mem['h1987] = 32'h206E776F;
mem['h1988] = 32'h6D6D6F63;
mem['h1989] = 32'h0D646E61;
mem['h198A] = 32'h0000000A;
mem['h198B] = 32'h00000000;
mem['h198C] = 32'h03020100;
mem['h198D] = 32'h07060504;
mem['h198E] = 32'h0B0A0908;
mem['h198F] = 32'h0F0E0D0C;
mem['h1990] = 32'h08040A0E;
mem['h1991] = 32'h060D0F09;
mem['h1992] = 32'h02000C01;
mem['h1993] = 32'h0305070B;
mem['h1994] = 32'h000C080B;
mem['h1995] = 32'h0D0F0205;
mem['h1996] = 32'h06030E0A;
mem['h1997] = 32'h04090107;
mem['h1998] = 32'h01030907;
mem['h1999] = 32'h0E0B0C0D;
mem['h199A] = 32'h0A050602;
mem['h199B] = 32'h080F0004;
mem['h199C] = 32'h07050009;
mem['h199D] = 32'h0F0A0402;
mem['h199E] = 32'h0C0B010E;
mem['h199F] = 32'h0D030806;
mem['h19A0] = 32'h0A060C02;
mem['h19A1] = 32'h03080B00;
mem['h19A2] = 32'h05070D04;
mem['h19A3] = 32'h09010E0F;
mem['h19A4] = 32'h0F01050C;
mem['h19A5] = 32'h0A040D0E;
mem['h19A6] = 32'h03060700;
mem['h19A7] = 32'h0B080209;
mem['h19A8] = 32'h0E070B0D;
mem['h19A9] = 32'h0903010C;
mem['h19AA] = 32'h040F0005;
mem['h19AB] = 32'h0A020608;
mem['h19AC] = 32'h090E0F06;
mem['h19AD] = 32'h0800030B;
mem['h19AE] = 32'h070D020C;
mem['h19AF] = 32'h050A0401;
mem['h19B0] = 32'h0408020A;
mem['h19B1] = 32'h05010607;
mem['h19B2] = 32'h0E090B0F;
mem['h19B3] = 32'h000D0C03;
mem['h19B4] = 32'h6A09E667;
mem['h19B5] = 32'hBB67AE85;
mem['h19B6] = 32'h3C6EF372;
mem['h19B7] = 32'hA54FF53A;
mem['h19B8] = 32'h510E527F;
mem['h19B9] = 32'h9B05688C;
mem['h19BA] = 32'h1F83D9AB;
mem['h19BB] = 32'h5BE0CD19;
mem['h19BC] = 32'h0000DB41;
mem['h19BD] = 32'h00000000;
mem['h19BE] = 32'h00000001;
mem['h19BF] = 32'h00000000;
mem['h19C0] = 32'h00000000;
mem['h19C1] = 32'h00000000;
mem['h19C2] = 32'h00000000;
mem['h19C3] = 32'h00000000;
mem['h19C4] = 32'h00000000;
mem['h19C5] = 32'h00000000;
mem['h19C6] = 32'h00000000;
mem['h19C7] = 32'h00000000;
mem['h19C8] = 32'h00000000;
mem['h19C9] = 32'h00000000;
mem['h19CA] = 32'h00000000;
mem['h19CB] = 32'h00000000;
mem['h19CC] = 32'h00000000;
mem['h19CD] = 32'h00000000;
mem['h19CE] = 32'h00000000;
mem['h19CF] = 32'h00000000;
mem['h19D0] = 32'h00000000;
mem['h19D1] = 32'h00000000;
mem['h19D2] = 32'h00000000;
mem['h19D3] = 32'h00000000;
mem['h19D4] = 32'h00000000;
mem['h19D5] = 32'h00000000;
mem['h19D6] = 32'h00000000;
mem['h19D7] = 32'h00000000;
mem['h19D8] = 32'h00000000;
mem['h19D9] = 32'h00000000;
mem['h19DA] = 32'h00000000;
mem['h19DB] = 32'h00000000;
mem['h19DC] = 32'h00000007;
mem['h19DD] = 32'h43424140;
mem['h19DE] = 32'h47464544;
mem['h19DF] = 32'h000059D4;
mem['h19E0] = 32'h307A2169;
mem['h19E1] = 32'h94809079;
mem['h19E2] = 32'hD02111E1;
mem['h19E3] = 32'h7C4A3542;
mem['h19E4] = 32'h48B6551F;
mem['h19E5] = 32'h1EA5A12C;
mem['h19E6] = 32'hFD0D251B;
mem['h19E7] = 32'hF9EED01E;
mem['h19E8] = 32'h00005BC0;
mem['h19E9] = 32'h8C5E8C50;
mem['h19EA] = 32'hE2147C32;
mem['h19EB] = 32'hA32BA7E1;
mem['h19EC] = 32'h2F45EB4E;
mem['h19ED] = 32'h208B4537;
mem['h19EE] = 32'h293AD69E;
mem['h19EF] = 32'h4C9B994D;
mem['h19F0] = 32'h82596786;
mem['h19F1] = 32'h00000009;
mem['h19F2] = 32'h00000000;
mem['h19F3] = 32'h00000000;
mem['h19F4] = 32'h00000000;
mem['h19F5] = 32'h00000000;
mem['h19F6] = 32'h00000000;
mem['h19F7] = 32'h00000000;
mem['h19F8] = 32'h00000000;
