-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
use work.global_wires_pkg.all;
-- Submodules: 975
entity tb_0CLK_447ec4ab is
port(
 clk : in std_logic;
 CLOCK_ENABLE : in unsigned(0 downto 0);
 global_to_module : in tb_global_to_module_t;
 module_to_global : out tb_module_to_global_t;
 return_output : out axis128_t_stream_t);
end tb_0CLK_447ec4ab;
architecture arch of tb_0CLK_447ec4ab is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function

-- All user state registers
signal input_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal ciphertext_in_stream : uint8_t_144 := (others => to_unsigned(0, 8));
signal ciphertext_remaining_in : unsigned(31 downto 0) := to_unsigned(0, 32);
signal cycle_counter : unsigned(31 downto 0) := to_unsigned(0, 32);
signal output_packet_count : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_size : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_remaining_out : unsigned(31 downto 0) := to_unsigned(0, 32);
signal plaintext_out_expected : char_128 := (others => to_unsigned(0, 8));
signal tag_match_checked : unsigned(0 downto 0) := to_unsigned(0, 1);
signal chacha20poly1305_decrypt_axis_in : axis128_t_stream_t := axis128_t_stream_t_NULL;
signal REG_COMB_input_packet_count : unsigned(31 downto 0);
signal REG_COMB_ciphertext_in_stream : uint8_t_144;
signal REG_COMB_ciphertext_remaining_in : unsigned(31 downto 0);
signal REG_COMB_cycle_counter : unsigned(31 downto 0);
signal REG_COMB_output_packet_count : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_size : unsigned(31 downto 0);
signal REG_COMB_plaintext_remaining_out : unsigned(31 downto 0);
signal REG_COMB_plaintext_out_expected : char_128;
signal REG_COMB_tag_match_checked : unsigned(0 downto 0);
signal REG_COMB_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;

-- Resolved maybe from input reg clock enable
signal clk_en_internal : std_logic;
-- Each function instance gets signals
-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l173_c8_1e61]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l174_c1_d93f]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output : unsigned(0 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(31 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : char_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : uint8_t_144;

-- printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7[chacha20poly1305_decrypt_tb_c_l175_c9_0af7]
signal printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_CLOCK_ENABLE : unsigned(0 downto 0);

-- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l177_c117_37e2]
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_x : unsigned(255 downto 0);
signal CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output : unsigned(255 downto 0);

-- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l177_c148_d32e]
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_x : unsigned(255 downto 0);
signal CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output : unsigned(255 downto 0);

-- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l177_c179_d9fe]
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_x : unsigned(255 downto 0);
signal CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output : unsigned(255 downto 0);

-- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l177_c210_7fa6]
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_x : unsigned(255 downto 0);
signal CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output : unsigned(255 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l177_c241_51ef]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_x : unsigned(255 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output : unsigned(255 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l177_c272_6b8d]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_x : unsigned(255 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output : unsigned(255 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l177_c302_2b93]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_x : unsigned(255 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output : unsigned(255 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l177_c332_b020]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_x : unsigned(255 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output : unsigned(255 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008[chacha20poly1305_decrypt_tb_c_l177_c64_3008]
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg3 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg4 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg5 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg6 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg7 : unsigned(31 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l178_c100_469b]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_x : unsigned(95 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output : unsigned(95 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l178_c130_1425]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_x : unsigned(95 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output : unsigned(95 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l178_c160_4e80]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_x : unsigned(95 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output : unsigned(95 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38[chacha20poly1305_decrypt_tb_c_l178_c65_8a38]
signal printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg2 : unsigned(31 downto 0);

-- print_aad[chacha20poly1305_decrypt_tb_c_l179_c9_781b]
signal print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_CLOCK_ENABLE : unsigned(0 downto 0);
signal print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad : uint8_t_32;
signal print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad_len : unsigned(31 downto 0);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l182_c32_f67f]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l183_c35_241b]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7[chacha20poly1305_decrypt_tb_c_l184_c9_05a7]
signal printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg1 : unsigned(31 downto 0);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l187_c30_1a07]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l190_c34_5523]
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_0 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_1 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output : char_array_128_t;

-- printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e[chacha20poly1305_decrypt_tb_c_l192_c9_5d0e]
signal printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l200_c8_abef]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_right : unsigned(0 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l201_c1_1f18]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(31 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(31 downto 0);

-- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : axis128_t_stream_t;
signal chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : axis128_t_stream_t;

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2]
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);

-- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l213_c56_ca58]
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_left : unsigned(31 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_right : unsigned(4 downto 0);
signal BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l216_c12_38ae]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l217_c1_0485]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(31 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(31 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l218_c176_9ef3]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l218_c207_36cf]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l218_c237_3380]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l218_c267_24cf]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25[chacha20poly1305_decrypt_tb_c_l218_c108_dc25]
signal printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg3 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l220_c1_ea25]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output : unsigned(0 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(31 downto 0);

-- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(31 downto 0);
signal input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(31 downto 0);

-- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef]
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
signal ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0[chacha20poly1305_decrypt_tb_c_l221_c17_56b0]
signal printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l223_c17_3079]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l225_c17_0ebd]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output : unsigned(31 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l234_c8_e9ad]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l235_c1_032c]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);

-- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l237_c169_597f]
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_x : unsigned(127 downto 0);
signal CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output : unsigned(127 downto 0);

-- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l237_c200_d957]
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_x : unsigned(127 downto 0);
signal CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output : unsigned(127 downto 0);

-- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l237_c230_8274]
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_x : unsigned(127 downto 0);
signal CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output : unsigned(127 downto 0);

-- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l237_c260_439a]
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_x : unsigned(127 downto 0);
signal CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output : unsigned(127 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77[chacha20poly1305_decrypt_tb_c_l237_c105_9a77]
signal printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg1 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg2 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg3 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951]
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
signal FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l254_c1_0e8a]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l261_c1_8ede]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l255_c16_51fa]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_right : unsigned(4 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l255_c1_a50b]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_a633]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l255_c13_ead1]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8[chacha20poly1305_decrypt_tb_c_l256_c17_35f8]
signal printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_CLOCK_ENABLE : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c[chacha20poly1305_decrypt_tb_c_l258_c17_2a1c]
signal printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_arg0 : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l262_c16_0389]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l262_c1_116d]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9]
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
signal plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96[chacha20poly1305_decrypt_tb_c_l263_c18_9c96]
signal printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_CLOCK_ENABLE : unsigned(0 downto 0);

-- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l265_c17_a77d]
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_right : unsigned(4 downto 0);
signal BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output : unsigned(31 downto 0);

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l272_c9_d81d]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_right : unsigned(0 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output : unsigned(0 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l272_c41_b474]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l272_c9_c63b]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output : unsigned(0 downto 0);

-- UNARY_OP_NOT[chacha20poly1305_decrypt_tb_c_l272_c69_ec38]
signal UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_expr : unsigned(0 downto 0);
signal UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output : unsigned(0 downto 0);

-- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l272_c9_dd50]
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_left : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_right : unsigned(0 downto 0);
signal BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l273_c1_c4e6]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output : unsigned(0 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(0 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);

-- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
signal output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : char_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : uint8_t_144;

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l275_c1_e50f]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output : unsigned(0 downto 0);

-- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l277_c1_ea4e]
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_cond : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iftrue : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iffalse : unsigned(0 downto 0);
signal FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output : unsigned(0 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7[chacha20poly1305_decrypt_tb_c_l276_c13_2af7]
signal printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_arg0 : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87[chacha20poly1305_decrypt_tb_c_l278_c13_ab87]
signal printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_arg0 : unsigned(31 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l282_c9_7928]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output : unsigned(32 downto 0);

-- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l283_c12_163a]
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_left : unsigned(31 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_right : unsigned(1 downto 0);
signal BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l284_c1_88f0]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output : unsigned(0 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : unsigned(31 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : char_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : uint8_t_144;

-- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l286_c17_1b46]
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_left : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_right : unsigned(31 downto 0);
signal BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output : unsigned(0 downto 0);

-- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l286_c1_c205]
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_cond : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iftrue : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iffalse : unsigned(0 downto 0);
signal TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output : unsigned(0 downto 0);

-- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea]
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : unsigned(31 downto 0);
signal plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : unsigned(31 downto 0);

-- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea]
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : unsigned(31 downto 0);
signal plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : unsigned(31 downto 0);

-- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea]
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : unsigned(31 downto 0);
signal ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : unsigned(31 downto 0);

-- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea]
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : char_128;
signal plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : char_128;

-- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea]
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : uint8_t_144;
signal ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : uint8_t_144;

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l288_c40_1f85]
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_0 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_1 : uint8_t_144;
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output : uint8_t_array_144_t;

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l289_c43_c7a8]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output : unsigned(31 downto 0);

-- printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec[chacha20poly1305_decrypt_tb_c_l290_c17_c7ec]
signal printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg1 : unsigned(31 downto 0);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l293_c38_2873]
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_0 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_1 : unsigned(31 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output : unsigned(31 downto 0);

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l296_c42_2383]
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_0 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_1 : char_128;
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_var_dim_0 : unsigned(0 downto 0);
signal VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output : char_array_128_t;

-- printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9[chacha20poly1305_decrypt_tb_c_l298_c17_cae9]
signal printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_CLOCK_ENABLE : unsigned(0 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg0 : unsigned(31 downto 0);
signal printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg1 : unsigned(31 downto 0);

-- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l305_c9_276d]
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_left : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_right : unsigned(31 downto 0);
signal BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output : unsigned(0 downto 0);

-- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l305_c5_427d]
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_cond : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iftrue : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iffalse : unsigned(0 downto 0);
signal tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output : unsigned(0 downto 0);

-- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l309_c5_c101]
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_left : unsigned(31 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_right : unsigned(0 downto 0);
signal BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output : unsigned(32 downto 0);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_left : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_right : unsigned(31 downto 0);
signal BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output : unsigned(31 downto 0);

function CONST_REF_RD_uint8_t_144_uint8_t_144_a26f( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_b938( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(0) := ref_toks_1;
      base(1) := ref_toks_2;
      base(2) := ref_toks_3;
      base(3) := ref_toks_4;
      base(4) := ref_toks_5;
      base(5) := ref_toks_6;
      base(6) := ref_toks_7;
      base(7) := ref_toks_8;
      base(8) := ref_toks_9;
      base(9) := ref_toks_10;
      base(10) := ref_toks_11;
      base(11) := ref_toks_12;
      base(12) := ref_toks_13;
      base(13) := ref_toks_14;
      base(14) := ref_toks_15;
      base(15) := ref_toks_16;
      base(16) := ref_toks_17;
      base(17) := ref_toks_18;
      base(18) := ref_toks_19;
      base(19) := ref_toks_20;
      base(20) := ref_toks_21;
      base(21) := ref_toks_22;
      base(22) := ref_toks_23;
      base(23) := ref_toks_24;
      base(24) := ref_toks_25;
      base(25) := ref_toks_26;
      base(26) := ref_toks_27;
      base(27) := ref_toks_28;
      base(28) := ref_toks_29;
      base(29) := ref_toks_30;
      base(30) := ref_toks_31;
      base(31) := ref_toks_32;
      base(32) := ref_toks_33;
      base(33) := ref_toks_34;
      base(34) := ref_toks_35;
      base(35) := ref_toks_36;
      base(36) := ref_toks_37;
      base(37) := ref_toks_38;
      base(38) := ref_toks_39;
      base(39) := ref_toks_40;
      base(40) := ref_toks_41;
      base(41) := ref_toks_42;
      base(42) := ref_toks_43;
      base(43) := ref_toks_44;
      base(44) := ref_toks_45;
      base(45) := ref_toks_46;
      base(46) := ref_toks_47;
      base(47) := ref_toks_48;
      base(48) := ref_toks_49;
      base(49) := ref_toks_50;
      base(50) := ref_toks_51;
      base(51) := ref_toks_52;
      base(52) := ref_toks_53;
      base(53) := ref_toks_54;
      base(54) := ref_toks_55;
      base(55) := ref_toks_56;
      base(56) := ref_toks_57;
      base(57) := ref_toks_58;
      base(58) := ref_toks_59;
      base(59) := ref_toks_60;
      base(60) := ref_toks_61;
      base(61) := ref_toks_62;
      base(62) := ref_toks_63;
      base(63) := ref_toks_64;
      base(64) := ref_toks_65;
      base(65) := ref_toks_66;
      base(66) := ref_toks_67;
      base(67) := ref_toks_68;
      base(68) := ref_toks_69;
      base(69) := ref_toks_70;
      base(70) := ref_toks_71;
      base(71) := ref_toks_72;
      base(72) := ref_toks_73;
      base(73) := ref_toks_74;
      base(74) := ref_toks_75;
      base(75) := ref_toks_76;
      base(76) := ref_toks_77;
      base(77) := ref_toks_78;
      base(78) := ref_toks_79;
      base(79) := ref_toks_80;
      base(80) := ref_toks_81;
      base(81) := ref_toks_82;
      base(82) := ref_toks_83;
      base(83) := ref_toks_84;
      base(84) := ref_toks_85;
      base(85) := ref_toks_86;
      base(86) := ref_toks_87;
      base(87) := ref_toks_88;
      base(88) := ref_toks_89;
      base(89) := ref_toks_90;
      base(90) := ref_toks_91;
      base(91) := ref_toks_92;
      base(92) := ref_toks_93;
      base(93) := ref_toks_94;
      base(94) := ref_toks_95;
      base(95) := ref_toks_96;

      return_output := base;
      return return_output; 
end function;

function uint8_array32_be( x : uint8_t_32) return unsigned is

  --variable x : uint8_t_32;
  variable return_output : unsigned(255 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15)&x(16)&x(17)&x(18)&x(19)&x(20)&x(21)&x(22)&x(23)&x(24)&x(25)&x(26)&x(27)&x(28)&x(29)&x(30)&x(31);
return return_output;
end function;

function uint8_array12_be( x : uint8_t_12) return unsigned is

  --variable x : uint8_t_12;
  variable return_output : unsigned(95 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11);
return return_output;
end function;

function CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned) return uint8_t_16 is
 
  variable base : axis128_t_stream_t; 
  variable return_output : uint8_t_16;
begin
      base.data.tdata(0) := ref_toks_0;
      base.data.tdata(1) := ref_toks_1;
      base.data.tdata(2) := ref_toks_2;
      base.data.tdata(3) := ref_toks_3;
      base.data.tdata(4) := ref_toks_4;
      base.data.tdata(5) := ref_toks_5;
      base.data.tdata(6) := ref_toks_6;
      base.data.tdata(7) := ref_toks_7;
      base.data.tdata(8) := ref_toks_8;
      base.data.tdata(9) := ref_toks_9;
      base.data.tdata(10) := ref_toks_10;
      base.data.tdata(11) := ref_toks_11;
      base.data.tdata(12) := ref_toks_12;
      base.data.tdata(13) := ref_toks_13;
      base.data.tdata(14) := ref_toks_14;
      base.data.tdata(15) := ref_toks_15;

      return_output := base.data.tdata;
      return return_output; 
end function;

function uint8_array16_be( x : uint8_t_16) return unsigned is

  --variable x : uint8_t_16;
  variable return_output : unsigned(127 downto 0);

begin
return_output := x(0)&x(1)&x(2)&x(3)&x(4)&x(5)&x(6)&x(7)&x(8)&x(9)&x(10)&x(11)&x(12)&x(13)&x(14)&x(15);
return return_output;
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base.data.tkeep(0) := ref_toks_0;
      base.data.tdata(0) := ref_toks_1;
      base.data.tkeep(1) := ref_toks_2;
      base.data.tdata(1) := ref_toks_3;
      base.data.tkeep(2) := ref_toks_4;
      base.data.tdata(2) := ref_toks_5;
      base.data.tkeep(3) := ref_toks_6;
      base.data.tdata(3) := ref_toks_7;
      base.data.tkeep(4) := ref_toks_8;
      base.data.tdata(4) := ref_toks_9;
      base.data.tkeep(5) := ref_toks_10;
      base.data.tdata(5) := ref_toks_11;
      base.data.tkeep(6) := ref_toks_12;
      base.data.tdata(6) := ref_toks_13;
      base.data.tkeep(7) := ref_toks_14;
      base.data.tdata(7) := ref_toks_15;
      base.data.tkeep(8) := ref_toks_16;
      base.data.tdata(8) := ref_toks_17;
      base.data.tkeep(9) := ref_toks_18;
      base.data.tdata(9) := ref_toks_19;
      base.data.tkeep(10) := ref_toks_20;
      base.data.tdata(10) := ref_toks_21;
      base.data.tkeep(11) := ref_toks_22;
      base.data.tdata(11) := ref_toks_23;
      base.data.tkeep(12) := ref_toks_24;
      base.data.tdata(12) := ref_toks_25;
      base.data.tkeep(13) := ref_toks_26;
      base.data.tdata(13) := ref_toks_27;
      base.data.tkeep(14) := ref_toks_28;
      base.data.tdata(14) := ref_toks_29;
      base.data.tkeep(15) := ref_toks_30;
      base.data.tdata(15) := ref_toks_31;
      base.data.tlast := ref_toks_32;
      base.valid := ref_toks_33;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee( ref_toks_0 : axis128_t_stream_t;
 ref_toks_1 : unsigned) return axis128_t_stream_t is
 
  variable base : axis128_t_stream_t; 
  variable return_output : axis128_t_stream_t;
begin
      base := ref_toks_0;
      base.valid := ref_toks_1;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_32_uint8_t_32_1367( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned) return uint8_t_32 is
 
  variable base : uint8_t_32; 
  variable return_output : uint8_t_32;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;
      base(12) := ref_toks_12;
      base(13) := ref_toks_13;
      base(14) := ref_toks_14;
      base(15) := ref_toks_15;
      base(16) := ref_toks_16;
      base(17) := ref_toks_17;
      base(18) := ref_toks_18;
      base(19) := ref_toks_19;
      base(20) := ref_toks_20;
      base(21) := ref_toks_21;
      base(22) := ref_toks_22;
      base(23) := ref_toks_23;
      base(24) := ref_toks_24;
      base(25) := ref_toks_25;
      base(26) := ref_toks_26;
      base(27) := ref_toks_27;
      base(28) := ref_toks_28;
      base(29) := ref_toks_29;
      base(30) := ref_toks_30;
      base(31) := ref_toks_31;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned) return uint8_t_12 is
 
  variable base : uint8_t_12; 
  variable return_output : uint8_t_12;
begin
      base(0) := ref_toks_0;
      base(1) := ref_toks_1;
      base(2) := ref_toks_2;
      base(3) := ref_toks_3;
      base(4) := ref_toks_4;
      base(5) := ref_toks_5;
      base(6) := ref_toks_6;
      base(7) := ref_toks_7;
      base(8) := ref_toks_8;
      base(9) := ref_toks_9;
      base(10) := ref_toks_10;
      base(11) := ref_toks_11;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_char_128_char_128_1091( ref_toks_0 : char_128;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned) return char_128 is
 
  variable base : char_128; 
  variable return_output : char_128;
begin
      base := ref_toks_0;
      base(108) := ref_toks_1;
      base(53) := ref_toks_2;
      base(50) := ref_toks_3;
      base(62) := ref_toks_4;
      base(59) := ref_toks_5;
      base(4) := ref_toks_6;
      base(68) := ref_toks_7;
      base(13) := ref_toks_8;
      base(77) := ref_toks_9;
      base(22) := ref_toks_10;
      base(19) := ref_toks_11;
      base(86) := ref_toks_12;
      base(83) := ref_toks_13;
      base(28) := ref_toks_14;
      base(92) := ref_toks_15;
      base(37) := ref_toks_16;
      base(101) := ref_toks_17;
      base(46) := ref_toks_18;
      base(110) := ref_toks_19;
      base(55) := ref_toks_20;
      base(52) := ref_toks_21;
      base(61) := ref_toks_22;
      base(6) := ref_toks_23;
      base(70) := ref_toks_24;
      base(15) := ref_toks_25;
      base(12) := ref_toks_26;
      base(79) := ref_toks_27;
      base(76) := ref_toks_28;
      base(21) := ref_toks_29;
      base(88) := ref_toks_30;
      base(85) := ref_toks_31;
      base(30) := ref_toks_32;
      base(94) := ref_toks_33;
      base(39) := ref_toks_34;
      base(103) := ref_toks_35;
      base(48) := ref_toks_36;
      base(45) := ref_toks_37;
      base(109) := ref_toks_38;
      base(54) := ref_toks_39;
      base(63) := ref_toks_40;
      base(8) := ref_toks_41;
      base(5) := ref_toks_42;
      base(72) := ref_toks_43;
      base(17) := ref_toks_44;
      base(69) := ref_toks_45;
      base(14) := ref_toks_46;
      base(81) := ref_toks_47;
      base(78) := ref_toks_48;
      base(23) := ref_toks_49;
      base(87) := ref_toks_50;
      base(32) := ref_toks_51;
      base(96) := ref_toks_52;
      base(41) := ref_toks_53;
      base(105) := ref_toks_54;
      base(38) := ref_toks_55;
      base(102) := ref_toks_56;
      base(47) := ref_toks_57;
      base(111) := ref_toks_58;
      base(56) := ref_toks_59;
      base(1) := ref_toks_60;
      base(65) := ref_toks_61;
      base(10) := ref_toks_62;
      base(7) := ref_toks_63;
      base(74) := ref_toks_64;
      base(71) := ref_toks_65;
      base(16) := ref_toks_66;
      base(80) := ref_toks_67;
      base(25) := ref_toks_68;
      base(89) := ref_toks_69;
      base(34) := ref_toks_70;
      base(98) := ref_toks_71;
      base(31) := ref_toks_72;
      base(43) := ref_toks_73;
      base(95) := ref_toks_74;
      base(107) := ref_toks_75;
      base(40) := ref_toks_76;
      base(104) := ref_toks_77;
      base(49) := ref_toks_78;
      base(58) := ref_toks_79;
      base(3) := ref_toks_80;
      base(0) := ref_toks_81;
      base(67) := ref_toks_82;
      base(64) := ref_toks_83;
      base(9) := ref_toks_84;
      base(73) := ref_toks_85;
      base(18) := ref_toks_86;
      base(82) := ref_toks_87;
      base(27) := ref_toks_88;
      base(91) := ref_toks_89;
      base(24) := ref_toks_90;
      base(36) := ref_toks_91;
      base(100) := ref_toks_92;
      base(33) := ref_toks_93;
      base(97) := ref_toks_94;
      base(42) := ref_toks_95;
      base(106) := ref_toks_96;
      base(51) := ref_toks_97;
      base(60) := ref_toks_98;
      base(57) := ref_toks_99;
      base(2) := ref_toks_100;
      base(66) := ref_toks_101;
      base(11) := ref_toks_102;
      base(75) := ref_toks_103;
      base(20) := ref_toks_104;
      base(84) := ref_toks_105;
      base(29) := ref_toks_106;
      base(93) := ref_toks_107;
      base(26) := ref_toks_108;
      base(90) := ref_toks_109;
      base(35) := ref_toks_110;
      base(99) := ref_toks_111;
      base(44) := ref_toks_112;

      return_output := base;
      return return_output; 
end function;

function CONST_REF_RD_uint8_t_144_uint8_t_144_10fa( ref_toks_0 : uint8_t_144;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned;
 ref_toks_5 : unsigned;
 ref_toks_6 : unsigned;
 ref_toks_7 : unsigned;
 ref_toks_8 : unsigned;
 ref_toks_9 : unsigned;
 ref_toks_10 : unsigned;
 ref_toks_11 : unsigned;
 ref_toks_12 : unsigned;
 ref_toks_13 : unsigned;
 ref_toks_14 : unsigned;
 ref_toks_15 : unsigned;
 ref_toks_16 : unsigned;
 ref_toks_17 : unsigned;
 ref_toks_18 : unsigned;
 ref_toks_19 : unsigned;
 ref_toks_20 : unsigned;
 ref_toks_21 : unsigned;
 ref_toks_22 : unsigned;
 ref_toks_23 : unsigned;
 ref_toks_24 : unsigned;
 ref_toks_25 : unsigned;
 ref_toks_26 : unsigned;
 ref_toks_27 : unsigned;
 ref_toks_28 : unsigned;
 ref_toks_29 : unsigned;
 ref_toks_30 : unsigned;
 ref_toks_31 : unsigned;
 ref_toks_32 : unsigned;
 ref_toks_33 : unsigned;
 ref_toks_34 : unsigned;
 ref_toks_35 : unsigned;
 ref_toks_36 : unsigned;
 ref_toks_37 : unsigned;
 ref_toks_38 : unsigned;
 ref_toks_39 : unsigned;
 ref_toks_40 : unsigned;
 ref_toks_41 : unsigned;
 ref_toks_42 : unsigned;
 ref_toks_43 : unsigned;
 ref_toks_44 : unsigned;
 ref_toks_45 : unsigned;
 ref_toks_46 : unsigned;
 ref_toks_47 : unsigned;
 ref_toks_48 : unsigned;
 ref_toks_49 : unsigned;
 ref_toks_50 : unsigned;
 ref_toks_51 : unsigned;
 ref_toks_52 : unsigned;
 ref_toks_53 : unsigned;
 ref_toks_54 : unsigned;
 ref_toks_55 : unsigned;
 ref_toks_56 : unsigned;
 ref_toks_57 : unsigned;
 ref_toks_58 : unsigned;
 ref_toks_59 : unsigned;
 ref_toks_60 : unsigned;
 ref_toks_61 : unsigned;
 ref_toks_62 : unsigned;
 ref_toks_63 : unsigned;
 ref_toks_64 : unsigned;
 ref_toks_65 : unsigned;
 ref_toks_66 : unsigned;
 ref_toks_67 : unsigned;
 ref_toks_68 : unsigned;
 ref_toks_69 : unsigned;
 ref_toks_70 : unsigned;
 ref_toks_71 : unsigned;
 ref_toks_72 : unsigned;
 ref_toks_73 : unsigned;
 ref_toks_74 : unsigned;
 ref_toks_75 : unsigned;
 ref_toks_76 : unsigned;
 ref_toks_77 : unsigned;
 ref_toks_78 : unsigned;
 ref_toks_79 : unsigned;
 ref_toks_80 : unsigned;
 ref_toks_81 : unsigned;
 ref_toks_82 : unsigned;
 ref_toks_83 : unsigned;
 ref_toks_84 : unsigned;
 ref_toks_85 : unsigned;
 ref_toks_86 : unsigned;
 ref_toks_87 : unsigned;
 ref_toks_88 : unsigned;
 ref_toks_89 : unsigned;
 ref_toks_90 : unsigned;
 ref_toks_91 : unsigned;
 ref_toks_92 : unsigned;
 ref_toks_93 : unsigned;
 ref_toks_94 : unsigned;
 ref_toks_95 : unsigned;
 ref_toks_96 : unsigned;
 ref_toks_97 : unsigned;
 ref_toks_98 : unsigned;
 ref_toks_99 : unsigned;
 ref_toks_100 : unsigned;
 ref_toks_101 : unsigned;
 ref_toks_102 : unsigned;
 ref_toks_103 : unsigned;
 ref_toks_104 : unsigned;
 ref_toks_105 : unsigned;
 ref_toks_106 : unsigned;
 ref_toks_107 : unsigned;
 ref_toks_108 : unsigned;
 ref_toks_109 : unsigned;
 ref_toks_110 : unsigned;
 ref_toks_111 : unsigned;
 ref_toks_112 : unsigned;
 ref_toks_113 : unsigned;
 ref_toks_114 : unsigned;
 ref_toks_115 : unsigned;
 ref_toks_116 : unsigned;
 ref_toks_117 : unsigned;
 ref_toks_118 : unsigned;
 ref_toks_119 : unsigned;
 ref_toks_120 : unsigned;
 ref_toks_121 : unsigned;
 ref_toks_122 : unsigned;
 ref_toks_123 : unsigned;
 ref_toks_124 : unsigned;
 ref_toks_125 : unsigned;
 ref_toks_126 : unsigned;
 ref_toks_127 : unsigned;
 ref_toks_128 : unsigned) return uint8_t_144 is
 
  variable base : uint8_t_144; 
  variable return_output : uint8_t_144;
begin
      base := ref_toks_0;
      base(100) := ref_toks_1;
      base(45) := ref_toks_2;
      base(109) := ref_toks_3;
      base(118) := ref_toks_4;
      base(11) := ref_toks_5;
      base(75) := ref_toks_6;
      base(20) := ref_toks_7;
      base(84) := ref_toks_8;
      base(29) := ref_toks_9;
      base(93) := ref_toks_10;
      base(38) := ref_toks_11;
      base(102) := ref_toks_12;
      base(47) := ref_toks_13;
      base(111) := ref_toks_14;
      base(4) := ref_toks_15;
      base(68) := ref_toks_16;
      base(13) := ref_toks_17;
      base(77) := ref_toks_18;
      base(22) := ref_toks_19;
      base(86) := ref_toks_20;
      base(31) := ref_toks_21;
      base(95) := ref_toks_22;
      base(40) := ref_toks_23;
      base(104) := ref_toks_24;
      base(61) := ref_toks_25;
      base(6) := ref_toks_26;
      base(125) := ref_toks_27;
      base(70) := ref_toks_28;
      base(15) := ref_toks_29;
      base(79) := ref_toks_30;
      base(24) := ref_toks_31;
      base(88) := ref_toks_32;
      base(33) := ref_toks_33;
      base(97) := ref_toks_34;
      base(54) := ref_toks_35;
      base(63) := ref_toks_36;
      base(8) := ref_toks_37;
      base(127) := ref_toks_38;
      base(72) := ref_toks_39;
      base(17) := ref_toks_40;
      base(81) := ref_toks_41;
      base(26) := ref_toks_42;
      base(90) := ref_toks_43;
      base(56) := ref_toks_44;
      base(1) := ref_toks_45;
      base(120) := ref_toks_46;
      base(65) := ref_toks_47;
      base(10) := ref_toks_48;
      base(74) := ref_toks_49;
      base(19) := ref_toks_50;
      base(83) := ref_toks_51;
      base(28) := ref_toks_52;
      base(92) := ref_toks_53;
      base(49) := ref_toks_54;
      base(113) := ref_toks_55;
      base(58) := ref_toks_56;
      base(3) := ref_toks_57;
      base(122) := ref_toks_58;
      base(67) := ref_toks_59;
      base(12) := ref_toks_60;
      base(76) := ref_toks_61;
      base(21) := ref_toks_62;
      base(85) := ref_toks_63;
      base(42) := ref_toks_64;
      base(106) := ref_toks_65;
      base(51) := ref_toks_66;
      base(115) := ref_toks_67;
      base(60) := ref_toks_68;
      base(5) := ref_toks_69;
      base(124) := ref_toks_70;
      base(69) := ref_toks_71;
      base(14) := ref_toks_72;
      base(78) := ref_toks_73;
      base(35) := ref_toks_74;
      base(99) := ref_toks_75;
      base(44) := ref_toks_76;
      base(108) := ref_toks_77;
      base(53) := ref_toks_78;
      base(117) := ref_toks_79;
      base(62) := ref_toks_80;
      base(7) := ref_toks_81;
      base(126) := ref_toks_82;
      base(71) := ref_toks_83;
      base(37) := ref_toks_84;
      base(101) := ref_toks_85;
      base(46) := ref_toks_86;
      base(110) := ref_toks_87;
      base(55) := ref_toks_88;
      base(0) := ref_toks_89;
      base(119) := ref_toks_90;
      base(64) := ref_toks_91;
      base(73) := ref_toks_92;
      base(30) := ref_toks_93;
      base(94) := ref_toks_94;
      base(39) := ref_toks_95;
      base(103) := ref_toks_96;
      base(48) := ref_toks_97;
      base(112) := ref_toks_98;
      base(57) := ref_toks_99;
      base(2) := ref_toks_100;
      base(121) := ref_toks_101;
      base(66) := ref_toks_102;
      base(23) := ref_toks_103;
      base(87) := ref_toks_104;
      base(32) := ref_toks_105;
      base(96) := ref_toks_106;
      base(41) := ref_toks_107;
      base(105) := ref_toks_108;
      base(50) := ref_toks_109;
      base(114) := ref_toks_110;
      base(59) := ref_toks_111;
      base(123) := ref_toks_112;
      base(16) := ref_toks_113;
      base(80) := ref_toks_114;
      base(25) := ref_toks_115;
      base(89) := ref_toks_116;
      base(34) := ref_toks_117;
      base(98) := ref_toks_118;
      base(43) := ref_toks_119;
      base(107) := ref_toks_120;
      base(52) := ref_toks_121;
      base(116) := ref_toks_122;
      base(9) := ref_toks_123;
      base(18) := ref_toks_124;
      base(82) := ref_toks_125;
      base(27) := ref_toks_126;
      base(91) := ref_toks_127;
      base(36) := ref_toks_128;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61 : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7 : entity work.printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_CLOCK_ENABLE);

-- CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2 : 0 clocks latency
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2 : entity work.CONST_SR_224_uint256_t_0CLK_de264c78 port map (
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_x,
CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output);

-- CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e : 0 clocks latency
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e : entity work.CONST_SR_192_uint256_t_0CLK_de264c78 port map (
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_x,
CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output);

-- CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe : 0 clocks latency
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe : entity work.CONST_SR_160_uint256_t_0CLK_de264c78 port map (
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_x,
CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output);

-- CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6 : 0 clocks latency
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6 : entity work.CONST_SR_128_uint256_t_0CLK_de264c78 port map (
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_x,
CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef : entity work.CONST_SR_96_uint256_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d : entity work.CONST_SR_64_uint256_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93 : entity work.CONST_SR_32_uint256_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020 : entity work.CONST_SR_0_uint256_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008 : entity work.printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg0,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg1,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg2,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg3,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg4,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg5,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg6,
printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg7);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b : entity work.CONST_SR_64_uint96_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425 : entity work.CONST_SR_32_uint96_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80 : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80 : entity work.CONST_SR_0_uint96_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38 : entity work.printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg0,
printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg1,
printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg2);

-- print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b : 0 clocks latency
print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b : entity work.print_aad_0CLK_fa355561 port map (
print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_CLOCK_ENABLE,
print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad,
print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad_len);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7 : entity work.printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg0,
printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg1);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output);

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523 : 0 clocks latency
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523 : entity work.VAR_REF_RD_char_128_char_2_128_VAR_90b8_0CLK_b45a16e1 port map (
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_1,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_var_dim_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e : entity work.printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg0,
printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef : entity work.BIN_OP_GT_uint32_t_uint1_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_axis128_t_stream_t_axis128_t_stream_t_0CLK_de264c78 port map (
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8 : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

-- BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58 : 0 clocks latency
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58 : entity work.BIN_OP_LTE_uint32_t_uint5_t_0CLK_e595f783 port map (
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_left,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_right,
BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0 : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3 : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3 : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380 : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25 : entity work.printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg0,
printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg1,
printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg2,
printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg3);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : 0 clocks latency
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef : entity work.MUX_uint1_t_uint8_t_uint8_t_0CLK_de264c78 port map (
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse,
ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0 : entity work.printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

-- CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f : 0 clocks latency
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f : entity work.CONST_SR_96_uint128_t_0CLK_de264c78 port map (
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_x,
CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output);

-- CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957 : 0 clocks latency
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957 : entity work.CONST_SR_64_uint128_t_0CLK_de264c78 port map (
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_x,
CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output);

-- CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274 : 0 clocks latency
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274 : entity work.CONST_SR_32_uint128_t_0CLK_de264c78 port map (
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_x,
CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output);

-- CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a : 0 clocks latency
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a : entity work.CONST_SR_0_uint128_t_0CLK_de264c78 port map (
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_x,
CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77 : entity work.printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg0,
printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg1,
printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg2,
printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg3);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a : entity work.BIN_OP_GT_int33_t_int32_t_0CLK_1aac2328 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200 : entity work.BIN_OP_NEQ_uint8_t_uint8_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882 : entity work.BIN_OP_PLUS_int33_t_int32_t_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output);

-- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : 0 clocks latency
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951 : entity work.printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_0CLK_de264c78 port map (
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1,
FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa : entity work.BIN_OP_GT_uint32_t_uint5_t_0CLK_5af1a430 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633 : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8 : entity work.printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_CLOCK_ENABLE);

-- printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c : entity work.printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_arg0);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389 : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : 0 clocks latency
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9 : entity work.MUX_uint1_t_char_char_0CLK_de264c78 port map (
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse,
plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96 : entity work.printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_CLOCK_ENABLE);

-- BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d : 0 clocks latency
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d : entity work.BIN_OP_MINUS_uint32_t_uint5_t_0CLK_de264c78 port map (
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_left,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_right,
BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d : entity work.BIN_OP_EQ_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474 : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474 : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output);

-- UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38 : 0 clocks latency
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38 : entity work.UNARY_OP_NOT_uint1_t_0CLK_de264c78 port map (
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_expr,
UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output);

-- BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50 : 0 clocks latency
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50 : entity work.BIN_OP_AND_uint1_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_left,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_right,
BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output);

-- FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e : 0 clocks latency
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_cond,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iftrue,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iffalse,
FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7 : entity work.printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_arg0);

-- printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87 : entity work.printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_arg0);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output);

-- BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a : 0 clocks latency
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a : entity work.BIN_OP_LT_uint32_t_uint2_t_0CLK_5af1a430 port map (
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_left,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_right,
BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2 : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output);

-- BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46 : 0 clocks latency
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46 : entity work.BIN_OP_EQ_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_left,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_right,
BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output);

-- TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205 : 0 clocks latency
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205 : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_cond,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iftrue,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iffalse,
TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output);

-- plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : 0 clocks latency
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse,
plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output);

-- plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : 0 clocks latency
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse,
plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output);

-- ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : 0 clocks latency
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse,
ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output);

-- plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : 0 clocks latency
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : entity work.MUX_uint1_t_char_128_char_128_0CLK_de264c78 port map (
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse,
plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output);

-- ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : 0 clocks latency
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea : entity work.MUX_uint1_t_uint8_t_144_uint8_t_144_0CLK_de264c78 port map (
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse,
ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output);

-- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85 : 0 clocks latency
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85 : entity work.VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_0CLK_e56a0f0b port map (
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_1,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_var_dim_0,
VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec : entity work.printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg0,
printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg1);

-- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873 : 0 clocks latency
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873 : entity work.VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_0CLK_9e8edf93 port map (
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_1,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_var_dim_0,
VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output);

-- VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383 : 0 clocks latency
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383 : entity work.VAR_REF_RD_char_128_char_2_128_VAR_90b8_0CLK_b45a16e1 port map (
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_1,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_var_dim_0,
VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output);

-- printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9 : 0 clocks latency
printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9 : entity work.printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_0CLK_de264c78 port map (
printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_CLOCK_ENABLE,
printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg0,
printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg1);

-- BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d : 0 clocks latency
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d : entity work.BIN_OP_GT_uint32_t_uint32_t_0CLK_380ecc95 port map (
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_left,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_right,
BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output);

-- tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d : 0 clocks latency
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_cond,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iftrue,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iffalse,
tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output);

-- BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101 : 0 clocks latency
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101 : entity work.BIN_OP_PLUS_uint32_t_uint1_t_0CLK_de264c78 port map (
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_left,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_right,
BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output);

-- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182 : 0 clocks latency
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182 : entity work.BIN_OP_MINUS_uint32_t_uint32_t_0CLK_de264c78 port map (
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_left,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_right,
BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output);



-- Resolve what clock enable to use for user logic
clk_en_internal <= CLOCK_ENABLE(0);
-- Combinatorial process for pipeline stages
process (
CLOCK_ENABLE,
clk_en_internal,
 -- Registers
 input_packet_count,
 ciphertext_in_stream,
 ciphertext_remaining_in,
 cycle_counter,
 output_packet_count,
 plaintext_out_size,
 plaintext_remaining_out,
 plaintext_out_expected,
 tag_match_checked,
 chacha20poly1305_decrypt_axis_in,
 -- Clock cross input
 global_to_module,
 -- All submodule outputs
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
 CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output,
 CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output,
 CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output,
 CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output,
 VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
 BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
 CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output,
 CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output,
 CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output,
 CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output,
 FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output,
 BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output,
 UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output,
 BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output,
 FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output,
 BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output,
 BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output,
 TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output,
 plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output,
 plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output,
 ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output,
 plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output,
 ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output,
 VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output,
 VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output,
 VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output,
 BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output,
 tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output,
 BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output,
 BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_key : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_nonce : uint8_t_12;
 variable VAR_chacha20poly1305_decrypt_aad : uint8_t_32;
 variable VAR_chacha20poly1305_decrypt_aad_len : unsigned(7 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out_ready : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_out : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_is_verified_out : unsigned(0 downto 0);
 variable VAR_key : uint8_t_32;
 variable VAR_nonce : uint8_t_12;
 variable VAR_aad : uint8_t_32;
 variable VAR_aad_len : unsigned(31 downto 0);
 variable VAR_aad_len_chacha20poly1305_decrypt_tb_c_l86_c14_5621_0 : unsigned(31 downto 0);
 variable VAR_plaintexts : char_2_128;
 variable VAR_plaintext_lens : uint32_t_2;
 variable VAR_input_ciphertext0 : uint8_t_144;
 variable VAR_input_ciphertext1 : uint8_t_144;
 variable VAR_input_ciphertexts : uint8_t_2_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l144_c9_f9bf_return_output : uint8_t_144;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l145_c9_1594_return_output : uint8_t_144;
 variable VAR_ciphertext_lens : uint32_t_2;
 variable VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l156_c5_57b8 : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : char_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l190_c9_e6e9 : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l182_c9_8fd6 : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_PRINT_32_BYTES_uint : unsigned(255 downto 0);
 variable VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg4 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg5 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg6 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_x : unsigned(255 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output : unsigned(255 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg7 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_x : unsigned(255 downto 0);
 variable VAR_PRINT_12_BYTES_uint : unsigned(95 downto 0);
 variable VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l178_c40_5e81_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_x : unsigned(95 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output : unsigned(95 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_x : unsigned(95 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad : uint8_t_32;
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad_len : unsigned(31 downto 0);
 variable VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output : char_array_128_t;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_0 : char_128;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_1 : char_128;
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : axis128_t_stream_t;
 variable VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond : unsigned(0 downto 0);
 variable VAR_i : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond : unsigned(0 downto 0);
 variable VAR_PRINT_16_BYTES_uint : unsigned(127 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l218_c62_4023_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l218_c45_791a_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_x : unsigned(127 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iffalse : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(31 downto 0);
 variable VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l223_c17_40d5 : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(31 downto 0);
 variable VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse : unsigned(7 downto 0);
 variable VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output : unsigned(31 downto 0);
 variable VAR_ARRAY_SHIFT_DOWN_i : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l234_c8_effa_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond : unsigned(0 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l237_c58_357d_return_output : uint8_t_16;
 variable VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l237_c41_5ef8_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg0 : unsigned(31 downto 0);
 variable VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg1 : unsigned(31 downto 0);
 variable VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_x : unsigned(127 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output : unsigned(127 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg3 : unsigned(31 downto 0);
 variable VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_x : unsigned(127 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_pos : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left : signed(32 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right : signed(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output : signed(33 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse : unsigned(7 downto 0);
 variable VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_right : unsigned(4 downto 0);
 variable VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output : unsigned(31 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_96_CONST_REF_RD_char_char_128_112_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_97_CONST_REF_RD_char_char_128_113_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_98_CONST_REF_RD_char_char_128_114_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_99_CONST_REF_RD_char_char_128_115_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_100_CONST_REF_RD_char_char_128_116_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_101_CONST_REF_RD_char_char_128_117_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_102_CONST_REF_RD_char_char_128_118_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_103_CONST_REF_RD_char_char_128_119_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_104_CONST_REF_RD_char_char_128_120_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_105_CONST_REF_RD_char_char_128_121_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_106_CONST_REF_RD_char_char_128_122_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_107_CONST_REF_RD_char_char_128_123_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_108_CONST_REF_RD_char_char_128_124_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_109_CONST_REF_RD_char_char_128_125_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_110_CONST_REF_RD_char_char_128_126_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_111_CONST_REF_RD_char_char_128_127_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_left : unsigned(0 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_left : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_expr : unsigned(0 downto 0);
 variable VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : unsigned(31 downto 0);
 variable VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451 : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : unsigned(31 downto 0);
 variable VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iffalse : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_cond : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iftrue : unsigned(0 downto 0);
 variable VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iffalse : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_arg0 : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output : unsigned(32 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_right : unsigned(1 downto 0);
 variable VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond : unsigned(0 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_cond : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iftrue : unsigned(0 downto 0);
 variable VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iffalse : unsigned(0 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : unsigned(31 downto 0);
 variable VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : unsigned(31 downto 0);
 variable VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : char_128;
 variable VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l296_c17_49ca : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : char_128;
 variable VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue : uint8_t_144;
 variable VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l288_c17_9f8c : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse : uint8_t_144;
 variable VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output : uint8_t_array_144_t;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_0 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_1 : uint8_t_144;
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_0 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_1 : unsigned(31 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_var_dim_0 : unsigned(0 downto 0);
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output : char_array_128_t;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_0 : char_128;
 variable VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_1 : char_128;
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg0 : unsigned(31 downto 0);
 variable VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg1 : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iftrue : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iffalse : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output : unsigned(0 downto 0);
 variable VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_cond : unsigned(0 downto 0);
 variable VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l309_c5_dcba : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_right : unsigned(0 downto 0);
 variable VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output : unsigned(32 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l153_l177_DUPLICATE_7f3f_return_output : uint8_t_32;
 variable VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l178_l154_DUPLICATE_dd41_return_output : uint8_t_12;
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_0f4e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output : unsigned(7 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_left : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_right : unsigned(31 downto 0);
 variable VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output : unsigned(31 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_8db9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_eef3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f7cb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_4ad9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_3f32_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f064_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_a1d4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_9de3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_fdc6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_fad4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_2b27_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_9afe_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_1e88_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_5650_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_dd23_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3_return_output : unsigned(7 downto 0);
 variable VAR_CONST_REF_RD_char_128_char_128_1091_chacha20poly1305_decrypt_tb_c_l283_l272_l286_DUPLICATE_d4fa_return_output : char_128;
 variable VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_10fa_chacha20poly1305_decrypt_tb_c_l286_l283_l272_DUPLICATE_f8a4_return_output : uint8_t_144;
 -- State registers comb logic variables
variable REG_VAR_input_packet_count : unsigned(31 downto 0);
variable REG_VAR_ciphertext_in_stream : uint8_t_144;
variable REG_VAR_ciphertext_remaining_in : unsigned(31 downto 0);
variable REG_VAR_cycle_counter : unsigned(31 downto 0);
variable REG_VAR_output_packet_count : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_size : unsigned(31 downto 0);
variable REG_VAR_plaintext_remaining_out : unsigned(31 downto 0);
variable REG_VAR_plaintext_out_expected : char_128;
variable REG_VAR_tag_match_checked : unsigned(0 downto 0);
variable REG_VAR_chacha20poly1305_decrypt_axis_in : axis128_t_stream_t;
begin

  -- STATE REGS
  -- Default read regs into vars
  REG_VAR_input_packet_count := input_packet_count;
  REG_VAR_ciphertext_in_stream := ciphertext_in_stream;
  REG_VAR_ciphertext_remaining_in := ciphertext_remaining_in;
  REG_VAR_cycle_counter := cycle_counter;
  REG_VAR_output_packet_count := output_packet_count;
  REG_VAR_plaintext_out_size := plaintext_out_size;
  REG_VAR_plaintext_remaining_out := plaintext_remaining_out;
  REG_VAR_plaintext_out_expected := plaintext_out_expected;
  REG_VAR_tag_match_checked := tag_match_checked;
  REG_VAR_chacha20poly1305_decrypt_axis_in := chacha20poly1305_decrypt_axis_in;
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(14, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(14, 32);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_right := to_unsigned(16, 5);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse := to_unsigned(0, 1);
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iffalse := to_unsigned(0, 32);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_1 := to_byte_array("PipelineC is the best HDL around :) Let's go CHILIChips Wireguard team!", 128);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(8, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(8, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(0, 32);
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_right := to_unsigned(16, 5);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(8, 32);
     VAR_aad_len_chacha20poly1305_decrypt_tb_c_l86_c14_5621_0 := to_unsigned(29, 32);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad_len := VAR_aad_len_chacha20poly1305_decrypt_tb_c_l86_c14_5621_0;
     VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l156_c5_57b8 := resize(VAR_aad_len_chacha20poly1305_decrypt_tb_c_l86_c14_5621_0, 8);
     VAR_chacha20poly1305_decrypt_aad_len := VAR_chacha20poly1305_decrypt_aad_len_chacha20poly1305_decrypt_tb_c_l156_c5_57b8;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_right := to_unsigned(1, 1);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_right := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iffalse := to_unsigned(0, 1);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iffalse := to_unsigned(0, 1);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_right := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(2, 32);
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_right := to_unsigned(16, 5);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(7, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(7, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_1 := to_unsigned(71, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_1 := to_unsigned(71, 32);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(10, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_0 := to_unsigned(56, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_0 := to_unsigned(56, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(15, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(15, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(10, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(15, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := to_unsigned(1, 1);
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_right := to_unsigned(1, 1);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_0 := to_byte_array("Hello CHILIChips - Wireguard team, let's test this aead!", 128);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iffalse := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(7, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_1 := to_unsigned(96, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_1 := to_unsigned(96, 32);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(13, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(13, 32);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_right := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(11, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(11, 32);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_right := to_unsigned(2, 2);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse := to_unsigned(0, 8);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(12, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(4, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(9, 32);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_right := to_unsigned(1, 1);
     VAR_chacha20poly1305_decrypt_axis_out_ready := to_unsigned(1, 1);
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_left := to_unsigned(1, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(1, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(1, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(1, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(9, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(14, 32);
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_right := to_unsigned(0, 1);
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_right := to_unsigned(2, 2);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(6, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(6, 32);
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iftrue := to_unsigned(0, 1);
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_right := to_unsigned(16, 5);
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iftrue := to_unsigned(0, 1);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iffalse := to_unsigned(0, 1);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(13, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_0 := to_unsigned(80, 32);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_0 := to_unsigned(80, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right := to_signed(5, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(2, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(2, 32);
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iffalse := to_unsigned(0, 1);
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad := to_byte_array("Additional authenticated data", 32);
     VAR_chacha20poly1305_decrypt_aad := to_byte_array("Additional authenticated data", 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := to_unsigned(0, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right := to_signed(3, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right := to_signed(3, 32);
     -- CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l153_l177_DUPLICATE_7f3f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l153_l177_DUPLICATE_7f3f_return_output := CONST_REF_RD_uint8_t_32_uint8_t_32_1367(
     to_unsigned(128, 8),
     to_unsigned(129, 8),
     to_unsigned(130, 8),
     to_unsigned(131, 8),
     to_unsigned(132, 8),
     to_unsigned(133, 8),
     to_unsigned(134, 8),
     to_unsigned(135, 8),
     to_unsigned(136, 8),
     to_unsigned(137, 8),
     to_unsigned(138, 8),
     to_unsigned(139, 8),
     to_unsigned(140, 8),
     to_unsigned(141, 8),
     to_unsigned(142, 8),
     to_unsigned(143, 8),
     to_unsigned(144, 8),
     to_unsigned(145, 8),
     to_unsigned(146, 8),
     to_unsigned(147, 8),
     to_unsigned(148, 8),
     to_unsigned(149, 8),
     to_unsigned(150, 8),
     to_unsigned(151, 8),
     to_unsigned(152, 8),
     to_unsigned(153, 8),
     to_unsigned(154, 8),
     to_unsigned(155, 8),
     to_unsigned(156, 8),
     to_unsigned(157, 8),
     to_unsigned(158, 8),
     to_unsigned(159, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_a26f[chacha20poly1305_decrypt_tb_c_l144_c9_f9bf] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l144_c9_f9bf_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_a26f(
     (others => to_unsigned(0, 8)),
     to_unsigned(215, 8),
     to_unsigned(30, 8),
     to_unsigned(133, 8),
     to_unsigned(49, 8),
     to_unsigned(110, 8),
     to_unsigned(221, 8),
     to_unsigned(3, 8),
     to_unsigned(242, 8),
     to_unsigned(92, 8),
     to_unsigned(174, 8),
     to_unsigned(198, 8),
     to_unsigned(184, 8),
     to_unsigned(94, 8),
     to_unsigned(232, 8),
     to_unsigned(122, 8),
     to_unsigned(221, 8),
     to_unsigned(225, 8),
     to_unsigned(237, 8),
     to_unsigned(168, 8),
     to_unsigned(104, 8),
     to_unsigned(96, 8),
     to_unsigned(115, 8),
     to_unsigned(11, 8),
     to_unsigned(185, 8),
     to_unsigned(168, 8),
     to_unsigned(235, 8),
     to_unsigned(162, 8),
     to_unsigned(227, 8),
     to_unsigned(117, 8),
     to_unsigned(246, 8),
     to_unsigned(102, 8),
     to_unsigned(196, 8),
     to_unsigned(35, 8),
     to_unsigned(178, 8),
     to_unsigned(235, 8),
     to_unsigned(84, 8),
     to_unsigned(201, 8),
     to_unsigned(250, 8),
     to_unsigned(121, 8),
     to_unsigned(88, 8),
     to_unsigned(152, 8),
     to_unsigned(174, 8),
     to_unsigned(215, 8),
     to_unsigned(124, 8),
     to_unsigned(142, 8),
     to_unsigned(251, 8),
     to_unsigned(38, 8),
     to_unsigned(128, 8),
     to_unsigned(28, 8),
     to_unsigned(119, 8),
     to_unsigned(146, 8),
     to_unsigned(15, 8),
     to_unsigned(219, 8),
     to_unsigned(8, 8),
     to_unsigned(9, 8),
     to_unsigned(110, 8),
     to_unsigned(96, 8),
     to_unsigned(164, 8),
     to_unsigned(133, 8),
     to_unsigned(207, 8),
     to_unsigned(17, 8),
     to_unsigned(184, 8),
     to_unsigned(27, 8),
     to_unsigned(89, 8),
     to_unsigned(93, 8),
     to_unsigned(168, 8),
     to_unsigned(125, 8),
     to_unsigned(106, 8),
     to_unsigned(45, 8),
     to_unsigned(3, 8),
     to_unsigned(201, 8),
     to_unsigned(186, 8),
     to_unsigned(223, 8),
     to_unsigned(92, 8),
     to_unsigned(185, 8),
     to_unsigned(71, 8),
     to_unsigned(116, 8),
     to_unsigned(66, 8),
     to_unsigned(18, 8),
     to_unsigned(63, 8));

     -- CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l178_l154_DUPLICATE_dd41 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l178_l154_DUPLICATE_dd41_return_output := CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2(
     to_unsigned(7, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(0, 8),
     to_unsigned(64, 8),
     to_unsigned(65, 8),
     to_unsigned(66, 8),
     to_unsigned(67, 8),
     to_unsigned(68, 8),
     to_unsigned(69, 8),
     to_unsigned(70, 8),
     to_unsigned(71, 8));

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_b938[chacha20poly1305_decrypt_tb_c_l145_c9_1594] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l145_c9_1594_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_b938(
     (others => to_unsigned(0, 8)),
     to_unsigned(207, 8),
     to_unsigned(18, 8),
     to_unsigned(153, 8),
     to_unsigned(56, 8),
     to_unsigned(109, 8),
     to_unsigned(148, 8),
     to_unsigned(46, 8),
     to_unsigned(223, 8),
     to_unsigned(86, 8),
     to_unsigned(194, 8),
     to_unsigned(230, 8),
     to_unsigned(136, 8),
     to_unsigned(22, 8),
     to_unsigned(245, 8),
     to_unsigned(98, 8),
     to_unsigned(203, 8),
     to_unsigned(225, 8),
     to_unsigned(162, 8),
     to_unsigned(237, 8),
     to_unsigned(76, 8),
     to_unsigned(125, 8),
     to_unsigned(33, 8),
     to_unsigned(38, 8),
     to_unsigned(154, 8),
     to_unsigned(145, 8),
     to_unsigned(170, 8),
     to_unsigned(177, 8),
     to_unsigned(245, 8),
     to_unsigned(58, 8),
     to_unsigned(247, 8),
     to_unsigned(109, 8),
     to_unsigned(193, 8),
     to_unsigned(110, 8),
     to_unsigned(164, 8),
     to_unsigned(226, 8),
     to_unsigned(24, 8),
     to_unsigned(224, 8),
     to_unsigned(235, 8),
     to_unsigned(42, 8),
     to_unsigned(12, 8),
     to_unsigned(203, 8),
     to_unsigned(250, 8),
     to_unsigned(213, 8),
     to_unsigned(96, 8),
     to_unsigned(218, 8),
     to_unsigned(152, 8),
     to_unsigned(26, 8),
     to_unsigned(161, 8),
     to_unsigned(57, 8),
     to_unsigned(77, 8),
     to_unsigned(241, 8),
     to_unsigned(6, 8),
     to_unsigned(215, 8),
     to_unsigned(25, 8),
     to_unsigned(30, 8),
     to_unsigned(111, 8),
     to_unsigned(55, 8),
     to_unsigned(205, 8),
     to_unsigned(247, 8),
     to_unsigned(170, 8),
     to_unsigned(118, 8),
     to_unsigned(205, 8),
     to_unsigned(122, 8),
     to_unsigned(43, 8),
     to_unsigned(152, 8),
     to_unsigned(145, 8),
     to_unsigned(176, 8),
     to_unsigned(58, 8),
     to_unsigned(35, 8),
     to_unsigned(116, 8),
     to_unsigned(207, 8),
     to_unsigned(172, 8),
     to_unsigned(236, 8),
     to_unsigned(106, 8),
     to_unsigned(222, 8),
     to_unsigned(195, 8),
     to_unsigned(78, 8),
     to_unsigned(102, 8),
     to_unsigned(105, 8),
     to_unsigned(120, 8),
     to_unsigned(7, 8),
     to_unsigned(199, 8),
     to_unsigned(227, 8),
     to_unsigned(31, 8),
     to_unsigned(15, 8),
     to_unsigned(235, 8),
     to_unsigned(75, 8),
     to_unsigned(97, 8),
     to_unsigned(234, 8),
     to_unsigned(45, 8),
     to_unsigned(210, 8),
     to_unsigned(164, 8),
     to_unsigned(89, 8),
     to_unsigned(124, 8),
     to_unsigned(174, 8),
     to_unsigned(233, 8));

     -- Submodule level 1
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l145_c9_1594_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_1 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_b938_chacha20poly1305_decrypt_tb_c_l145_c9_1594_return_output;
     VAR_chacha20poly1305_decrypt_nonce := VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l178_l154_DUPLICATE_dd41_return_output;
     VAR_chacha20poly1305_decrypt_key := VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l153_l177_DUPLICATE_7f3f_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l144_c9_f9bf_return_output;
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_0 := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_a26f_chacha20poly1305_decrypt_tb_c_l144_c9_f9bf_return_output;
     -- uint8_array12_be[chacha20poly1305_decrypt_tb_c_l178_c40_5e81] LATENCY=0
     VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l178_c40_5e81_return_output := uint8_array12_be(
     VAR_CONST_REF_RD_uint8_t_12_uint8_t_12_b0e2_chacha20poly1305_decrypt_tb_c_l178_l154_DUPLICATE_dd41_return_output);

     -- uint8_array32_be[chacha20poly1305_decrypt_tb_c_l177_c41_8eed] LATENCY=0
     VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output := uint8_array32_be(
     VAR_CONST_REF_RD_uint8_t_32_uint8_t_32_1367_chacha20poly1305_decrypt_tb_c_l153_l177_DUPLICATE_7f3f_return_output);

     -- Submodule level 2
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_x := VAR_uint8_array32_be_chacha20poly1305_decrypt_tb_c_l177_c41_8eed_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l178_c40_5e81_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l178_c40_5e81_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_x := VAR_uint8_array12_be_chacha20poly1305_decrypt_tb_c_l178_c40_5e81_return_output;
     -- CONST_SR_160[chacha20poly1305_decrypt_tb_c_l177_c179_d9fe] LATENCY=0
     -- Inputs
     CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_x <= VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_x;
     -- Outputs
     VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output := CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output;

     -- CONST_SR_128[chacha20poly1305_decrypt_tb_c_l177_c210_7fa6] LATENCY=0
     -- Inputs
     CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_x <= VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_x;
     -- Outputs
     VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output := CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l178_c130_1425] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l178_c160_4e80] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output;

     -- CONST_SR_192[chacha20poly1305_decrypt_tb_c_l177_c148_d32e] LATENCY=0
     -- Inputs
     CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_x <= VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_x;
     -- Outputs
     VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output := CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output;

     -- CONST_SR_224[chacha20poly1305_decrypt_tb_c_l177_c117_37e2] LATENCY=0
     -- Inputs
     CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_x <= VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_x;
     -- Outputs
     VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output := CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l178_c100_469b] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l177_c302_2b93] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l177_c241_51ef] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l177_c272_6b8d] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l177_c332_b020] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg3 := resize(VAR_CONST_SR_128_chacha20poly1305_decrypt_tb_c_l177_c210_7fa6_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg2 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l178_c160_4e80_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg0 := resize(VAR_CONST_SR_224_chacha20poly1305_decrypt_tb_c_l177_c117_37e2_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg7 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l177_c332_b020_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg2 := resize(VAR_CONST_SR_160_chacha20poly1305_decrypt_tb_c_l177_c179_d9fe_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg4 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l177_c241_51ef_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg0 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l178_c100_469b_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg6 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l177_c302_2b93_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg5 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l177_c272_6b8d_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg1 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l178_c130_1425_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg1 := resize(VAR_CONST_SR_192_chacha20poly1305_decrypt_tb_c_l177_c148_d32e_return_output, 32);
 -- Reads from global variables
     VAR_chacha20poly1305_decrypt_axis_in_ready := global_to_module.chacha20poly1305_decrypt_axis_in_ready;
     VAR_chacha20poly1305_decrypt_axis_out := global_to_module.chacha20poly1305_decrypt_axis_out;
     VAR_chacha20poly1305_decrypt_is_verified_out := global_to_module.chacha20poly1305_decrypt_is_verified_out;
     -- Submodule level 0
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_right := VAR_chacha20poly1305_decrypt_axis_in_ready;
     VAR_return_output := VAR_chacha20poly1305_decrypt_axis_out;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_cond := VAR_chacha20poly1305_decrypt_is_verified_out;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_cond := VAR_chacha20poly1305_decrypt_is_verified_out;
     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d[chacha20poly1305_decrypt_tb_c_l254_c12_8420] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tlast;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_a1d4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_a1d4_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(7);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_4ad9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_4ad9_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(4);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_1e88 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_1e88_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(13);

     -- CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d[chacha20poly1305_decrypt_tb_c_l234_c8_effa] LATENCY=0
     VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l234_c8_effa_return_output := VAR_chacha20poly1305_decrypt_axis_out.valid;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_eef3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_eef3_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(2);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_9de3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_9de3_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(8);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_5650 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_5650_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(14);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_9afe LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_9afe_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(12);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_2b27 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_2b27_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(11);

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d[chacha20poly1305_decrypt_tb_c_l237_c58_357d] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l237_c58_357d_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata;

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f064 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f064_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(6);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_fdc6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_fdc6_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(9);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_fad4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_fad4_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(10);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f7cb LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f7cb_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(3);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_0f4e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_0f4e_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(0);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_dd23 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_dd23_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(15);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_3f32 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_3f32_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(5);

     -- CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_8db9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_8db9_return_output := VAR_chacha20poly1305_decrypt_axis_out.data.tdata(1);

     -- Submodule level 1
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_a1d4_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_7_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_a1d4_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_left := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_valid_d41d_chacha20poly1305_decrypt_tb_c_l234_c8_effa_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_5650_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_5650_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_dd23_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_15_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_dd23_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f064_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_6_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f064_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_1e88_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_13_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_1e88_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_9de3_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_8_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_9de3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_fdc6_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_9_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_fdc6_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_9afe_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_12_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_9afe_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_fad4_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_10_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_fad4_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_3f32_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_3f32_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_8db9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_8db9_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_2b27_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_11_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_2b27_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f7cb_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_3_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_f7cb_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_0f4e_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_0_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_0f4e_return_output, 32);
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond := VAR_CONST_REF_RD_uint1_t_axis128_t_stream_t_data_tlast_d41d_chacha20poly1305_decrypt_tb_c_l254_c12_8420_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_eef3_return_output, 32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_2_d41d_chacha20poly1305_decrypt_tb_c_l248_l244_DUPLICATE_eef3_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left := VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_4ad9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 := resize(VAR_CONST_REF_RD_uint8_t_axis128_t_stream_t_data_tdata_4_d41d_chacha20poly1305_decrypt_tb_c_l244_l248_DUPLICATE_4ad9_return_output, 32);
     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l237_c41_5ef8] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l237_c41_5ef8_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_d41d_chacha20poly1305_decrypt_tb_c_l237_c58_357d_return_output);

     -- Submodule level 2
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l237_c41_5ef8_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l237_c41_5ef8_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l237_c41_5ef8_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l237_c41_5ef8_return_output;
     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l237_c200_d957] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l237_c169_597f] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l237_c230_8274] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output;

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l237_c260_439a] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output;

     -- Submodule level 3
     VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l237_c169_597f_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l237_c260_439a_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l237_c230_8274_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l237_c200_d957_return_output, 32);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in clock enable
     VAR_CLOCK_ENABLE(0) := clk_en_internal;

     -- Submodule level 0
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iftrue := VAR_CLOCK_ENABLE;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iftrue := VAR_CLOCK_ENABLE;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse := ciphertext_in_stream;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse := ciphertext_remaining_in;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_left := cycle_counter;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_left := input_packet_count;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_var_dim_0 := resize(input_packet_count, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_var_dim_0 := resize(input_packet_count, 1);
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := input_packet_count;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg0 := input_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_arg0 := input_packet_count;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_left := output_packet_count;
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_left := output_packet_count;
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_var_dim_0 := resize(output_packet_count, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_var_dim_0 := resize(output_packet_count, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_arg0 := output_packet_count;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_arg0 := output_packet_count;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse := plaintext_out_expected;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse := plaintext_out_size;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse := plaintext_remaining_out;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse := tag_match_checked;
     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l182_c32_f67f] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l183_c35_241b] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output;

     -- chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee(
     chacha20poly1305_decrypt_axis_in,
     to_unsigned(0, 1));

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l223_c17_3079] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l234_c8_e9ad] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l216_c12_38ae] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l282_c9_7928] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l187_c30_1a07] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l173_c8_1e61] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l272_c41_b474] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output;

     -- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l190_c34_5523] LATENCY=0
     -- Inputs
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_0;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_1 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_ref_toks_1;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_var_dim_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output := VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output;

     -- BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l309_c5_c101] LATENCY=0
     -- Inputs
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_left <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_left;
     BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_right <= VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_right;
     -- Outputs
     VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output := BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output;

     -- Submodule level 1
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l216_c12_38ae_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l234_c8_e9ad_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l173_c8_1e61_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_right := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l272_c41_b474_return_output;
     VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l223_c17_40d5 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l223_c17_3079_return_output, 32);
     VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451 := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l282_c9_7928_return_output, 32);
     VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l309_c5_dcba := resize(VAR_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l309_c5_c101_return_output, 32);
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l190_c9_e6e9 := VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l190_c34_5523_return_output.data;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l183_c35_241b_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l187_c30_1a07_return_output;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l182_c9_8fd6 := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l182_c32_f67f_return_output.data;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_chacha20poly1305_decrypt_axis_in_FALSE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_2dee_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l182_c9_8fd6;
     REG_VAR_cycle_counter := VAR_cycle_counter_chacha20poly1305_decrypt_tb_c_l309_c5_dcba;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_input_packet_count_chacha20poly1305_decrypt_tb_c_l223_c17_40d5;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_right := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451;
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_left := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451;
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451, 1);
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_var_dim_0 := resize(VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451, 1);
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg0 := VAR_output_packet_count_chacha20poly1305_decrypt_tb_c_l282_c9_c451;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l190_c9_e6e9;
     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l293_c38_2873] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l174_c1_d93f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;

     -- BIN_OP_LT[chacha20poly1305_decrypt_tb_c_l283_c12_163a] LATENCY=0
     -- Inputs
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_left <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_left;
     BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_right <= VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_right;
     -- Outputs
     VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output := BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l235_c1_032c] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;

     -- VAR_REF_RD_char_128_char_2_128_VAR_90b8[chacha20poly1305_decrypt_tb_c_l296_c42_2383] LATENCY=0
     -- Inputs
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_0;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_1 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_ref_toks_1;
     VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_var_dim_0 <= VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output := VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l173_c5_dd91] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;

     -- Submodule level 2
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond := VAR_BIN_OP_LT_chacha20poly1305_decrypt_tb_c_l283_c12_163a_return_output;
     VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l174_c1_d93f_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l235_c1_032c_return_output;
     VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l296_c17_49ca := VAR_VAR_REF_RD_char_128_char_2_128_VAR_90b8_chacha20poly1305_decrypt_tb_c_l296_c42_2383_return_output.data;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l293_c38_2873_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_left := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left := signed(std_logic_vector(resize(VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_left := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_right := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left := signed(std_logic_vector(resize(VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output, 33)));
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_expr := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue := VAR_plaintext_out_expected_chacha20poly1305_decrypt_tb_c_l296_c17_49ca;
     -- CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(53);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(139);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(106);

     -- CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(68);

     -- CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb LATENCY=0
     VAR_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(26);

     -- CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(120);

     -- CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(99);

     -- CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(54);

     -- CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(85);

     -- CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(17);

     -- CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(21);

     -- CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(81);

     -- CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(33);

     -- CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(60);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_106_CONST_REF_RD_char_char_128_122_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_106_CONST_REF_RD_char_char_128_122_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(122);

     -- CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d LATENCY=0
     VAR_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(20);

     -- CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(61);

     -- CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(106);

     -- CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(117);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(138);

     -- UNARY_OP_NOT[chacha20poly1305_decrypt_tb_c_l272_c69_ec38] LATENCY=0
     -- Inputs
     UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_expr <= VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_expr;
     -- Outputs
     VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output := UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(122);

     -- CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(48);

     -- CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(71);

     -- CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(34);

     -- CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(54);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l265_c17_a77d] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output;

     -- CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(75);

     -- CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(40);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77[chacha20poly1305_decrypt_tb_c_l237_c105_9a77] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_chacha20poly1305_decrypt_tb_c_l237_c105_9a77_arg3;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(57);

     -- printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38[chacha20poly1305_decrypt_tb_c_l178_c65_8a38] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_chacha20poly1305_decrypt_tb_c_l178_c65_8a38_arg2;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(16);

     -- CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef LATENCY=0
     VAR_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(69);

     -- CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(78);

     -- CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(89);

     -- CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(45);

     -- CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(40);

     -- printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008[chacha20poly1305_decrypt_tb_c_l177_c64_3008] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg3;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg4 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg4;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg5 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg5;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg6 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg6;
     printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg7 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l177_c64_3008_chacha20poly1305_decrypt_tb_c_l177_c64_3008_arg7;
     -- Outputs

     -- CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d LATENCY=0
     VAR_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(74);

     -- CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(107);

     -- CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(11);

     -- CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(66);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(134);

     -- CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(75);

     -- CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(31);

     -- CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(13);

     -- CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(92);

     -- CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(82);

     -- CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(0);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f LATENCY=0
     VAR_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(102);

     -- CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(96);

     -- CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(113);

     -- CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(110);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(137);

     -- CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(10);

     -- CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(51);

     -- CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(98);

     -- CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(53);

     -- CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a LATENCY=0
     VAR_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(19);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_105_CONST_REF_RD_char_char_128_121_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_105_CONST_REF_RD_char_char_128_121_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(121);

     -- CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(15);

     -- CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae LATENCY=0
     VAR_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(27);

     -- CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(11);

     -- CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(74);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_107_CONST_REF_RD_char_char_128_123_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_107_CONST_REF_RD_char_char_128_123_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(123);

     -- CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(50);

     -- CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(110);

     -- CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(49);

     -- CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(34);

     -- CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(39);

     -- printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7[chacha20poly1305_decrypt_tb_c_l175_c9_0af7] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_chacha20poly1305_decrypt_tb_c_l175_c9_0af7_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec LATENCY=0
     VAR_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(68);

     -- CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(55);

     -- CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(88);

     -- CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(35);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_100_CONST_REF_RD_char_char_128_116_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_100_CONST_REF_RD_char_char_128_116_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(116);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(136);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(83);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(44);

     -- CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(85);

     -- CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e LATENCY=0
     VAR_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(71);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(77);

     -- CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(109);

     -- CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(76);

     -- CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(4);

     -- CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(62);

     -- CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(127);

     -- CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(16);

     -- CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(63);

     -- CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(37);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(51);

     -- CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(22);

     -- CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(50);

     -- CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(82);

     -- CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(23);

     -- CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(108);

     -- CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(88);

     -- CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(100);

     -- CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(30);

     -- CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e LATENCY=0
     VAR_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(87);

     -- CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(108);

     -- CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(55);

     -- CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(86);

     -- CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(98);

     -- BIN_OP_LTE[chacha20poly1305_decrypt_tb_c_l213_c56_ca58] LATENCY=0
     -- Inputs
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_left <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_left;
     BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_right <= VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_right;
     -- Outputs
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output := BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;

     -- CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(95);

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l261_c1_8ede] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(31);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(79);

     -- CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(9);

     -- CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a LATENCY=0
     VAR_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(105);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(56);

     -- CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(32);

     -- CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(96);

     -- CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(60);

     -- CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(35);

     -- CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(20);

     -- CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(70);

     -- CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(14);

     -- CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(15);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(42);

     -- CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(27);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(67);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(47);

     -- CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(104);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b LATENCY=0
     VAR_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(73);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_103_CONST_REF_RD_char_char_128_119_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_103_CONST_REF_RD_char_char_128_119_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(119);

     -- CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(111);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(133);

     -- CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada LATENCY=0
     VAR_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(65);

     -- CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(32);

     -- CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(10);

     -- CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(112);

     -- CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(8);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(129);

     -- print_aad[chacha20poly1305_decrypt_tb_c_l179_c9_781b] LATENCY=0
     -- Clock enable
     print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_CLOCK_ENABLE <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_CLOCK_ENABLE;
     -- Inputs
     print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad;
     print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad_len <= VAR_print_aad_chacha20poly1305_decrypt_tb_c_l179_c9_781b_aad_len;
     -- Outputs

     -- CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc LATENCY=0
     VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(0);

     -- CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(43);

     -- CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac LATENCY=0
     VAR_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(22);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(58);

     -- CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(63);

     -- BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182 LATENCY=0
     -- Inputs
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_left <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_left;
     BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_right <= VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_right;
     -- Outputs
     VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output := BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(2);

     -- CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(76);

     -- CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(3);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_108_CONST_REF_RD_char_char_128_124_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_108_CONST_REF_RD_char_char_128_124_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(124);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_104_CONST_REF_RD_char_char_128_120_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_104_CONST_REF_RD_char_char_128_120_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(120);

     -- CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(21);

     -- CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(94);

     -- CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e LATENCY=0
     VAR_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(83);

     -- CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(45);

     -- CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(92);

     -- CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(6);

     -- CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(123);

     -- CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(116);

     -- CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(103);

     -- CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(13);

     -- CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(65);

     -- CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(95);

     -- CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(41);

     -- CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(19);

     -- CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(42);

     -- CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(47);

     -- CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(87);

     -- CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(90);

     -- CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac LATENCY=0
     VAR_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(80);

     -- CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa LATENCY=0
     VAR_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(99);

     -- CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(59);

     -- CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(57);

     -- CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(25);

     -- CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(38);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_98_CONST_REF_RD_char_char_128_114_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_98_CONST_REF_RD_char_char_128_114_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(114);

     -- CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(41);

     -- CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(52);

     -- CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(90);

     -- CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(62);

     -- CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd LATENCY=0
     VAR_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(18);

     -- CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(91);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(141);

     -- CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(36);

     -- CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb LATENCY=0
     VAR_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(39);

     -- CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(89);

     -- CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(28);

     -- CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf LATENCY=0
     VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(7);

     -- CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f LATENCY=0
     VAR_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(23);

     -- CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(6);

     -- CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(8);

     -- CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(38);

     -- CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(73);

     -- CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(64);

     -- CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(125);

     -- CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed LATENCY=0
     VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(3);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_101_CONST_REF_RD_char_char_128_117_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_101_CONST_REF_RD_char_char_128_117_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(117);

     -- CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(44);

     -- CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(29);

     -- CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(78);

     -- CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f LATENCY=0
     VAR_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(72);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(102);

     -- printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e[chacha20poly1305_decrypt_tb_c_l192_c9_5d0e] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_chacha20poly1305_decrypt_tb_c_l192_c9_5d0e_arg1;
     -- Outputs

     -- CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(84);

     -- CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(36);

     -- CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(101);

     -- CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(46);

     -- CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(93);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(130);

     -- CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(91);

     -- CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(58);

     -- CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(33);

     -- CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(86);

     -- CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(59);

     -- CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(25);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_110_CONST_REF_RD_char_char_128_126_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_110_CONST_REF_RD_char_char_128_126_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(126);

     -- CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(103);

     -- CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(24);

     -- CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(119);

     -- CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(111);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba LATENCY=0
     VAR_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(66);

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l254_c1_0e8a] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(115);

     -- CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(97);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(143);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(121);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l200_c8_abef] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;

     -- CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(43);

     -- CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(124);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_96_CONST_REF_RD_char_char_128_112_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_96_CONST_REF_RD_char_char_128_112_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(112);

     -- CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(94);

     -- CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f LATENCY=0
     VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(4);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(5);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(132);

     -- CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(49);

     -- CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(5);

     -- CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(28);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_99_CONST_REF_RD_char_char_128_115_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_99_CONST_REF_RD_char_char_128_115_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(115);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(142);

     -- CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(67);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_97_CONST_REF_RD_char_char_128_113_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_97_CONST_REF_RD_char_char_128_113_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(113);

     -- CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(7);

     -- CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(81);

     -- CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a LATENCY=0
     VAR_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(61);

     -- CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(118);

     -- CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(26);

     -- CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(24);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(128);

     -- CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(12);

     -- CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f LATENCY=0
     VAR_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(93);

     -- CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(79);

     -- CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(126);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(131);

     -- printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7[chacha20poly1305_decrypt_tb_c_l184_c9_05a7] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_chacha20poly1305_decrypt_tb_c_l184_c9_05a7_arg1;
     -- Outputs

     -- CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a LATENCY=0
     VAR_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(64);

     -- CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(70);

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l255_c16_51fa] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output;

     -- CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(9);

     -- CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(14);

     -- CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b LATENCY=0
     VAR_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(77);

     -- CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(12);

     -- CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(52);

     -- CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(1);

     -- CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(105);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(18);

     -- CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd LATENCY=0
     VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(1);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_111_CONST_REF_RD_char_char_128_127_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_111_CONST_REF_RD_char_char_128_127_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(127);

     -- CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(72);

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l262_c16_0389] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_109_CONST_REF_RD_char_char_128_125_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_109_CONST_REF_RD_char_char_128_125_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(125);

     -- CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(29);

     -- FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_102_CONST_REF_RD_char_char_128_118_d41d[chacha20poly1305_decrypt_tb_c_l266_c168_d9f8] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_102_CONST_REF_RD_char_char_128_118_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(118);

     -- CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(48);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(100);

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l207_c16_98a8] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_left;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;

     -- CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(104);

     -- CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(84);

     -- CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(109);

     -- CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(114);

     -- CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(30);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l242_c16_321a] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(135);

     -- CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c LATENCY=0
     VAR_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(107);

     -- CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(80);

     -- CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(56);

     -- CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc LATENCY=0
     VAR_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(37);

     -- FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d[chacha20poly1305_decrypt_tb_c_l226_c173_b5dd] LATENCY=0
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(140);

     -- CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(101);

     -- CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(46);

     -- CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc LATENCY=0
     VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc_return_output := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(69);

     -- CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(97);

     -- CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(17);

     -- BIN_OP_MINUS[chacha20poly1305_decrypt_tb_c_l225_c17_0ebd] LATENCY=0
     -- Inputs
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_left <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_left;
     BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_right <= VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_right;
     -- Outputs
     VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output := BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output;

     -- CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8 LATENCY=0
     VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output(2);

     -- Submodule level 3
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l262_c16_0389_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l200_c8_abef_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l255_c16_51fa_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond := VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l225_c17_0ebd_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_BIN_OP_MINUS_chacha20poly1305_decrypt_tb_c_l265_c17_a77d_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left := signed(std_logic_vector(resize(VAR_BIN_OP_MINUS_uint32_t_uint32_t_chacha20poly1305_decrypt_tb_c_l246_DUPLICATE_c182_return_output, 33)));
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output, 32);
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_0_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l262_l244_DUPLICATE_95dc_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_100_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_f97c_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_101_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_cb38_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_102_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_4e4f_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_103_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2db7_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_104_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_ab10_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_105_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_b81a_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_106_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_2606_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_107_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_307c_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_108_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_f7c9_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_109_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6cb7_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output, 32);
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_10_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l248_l262_l244_DUPLICATE_c322_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_110_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b2b9_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_111_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_5182_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output, 32);
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_11_d41d_chacha20poly1305_decrypt_tb_c_l262_l244_l234_l254_l248_DUPLICATE_bfb9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output, 32);
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_12_d41d_chacha20poly1305_decrypt_tb_c_l262_l248_l234_l254_l244_DUPLICATE_e1a0_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output, 32);
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_13_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l234_l254_l248_DUPLICATE_aa19_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output, 32);
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_14_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l254_l234_DUPLICATE_e138_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output, 32);
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_15_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l248_l244_DUPLICATE_eca1_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_16_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_eaa9_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_17_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_c607_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_18_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_b3fd_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_19_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_957a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output, 32);
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_1_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l254_l248_l234_DUPLICATE_9dbd_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_20_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_411d_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_21_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_5291_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_22_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_c6ac_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_23_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_5d6f_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_24_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_17a3_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_25_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_0398_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_26_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_2abb_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_27_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l266_l234_DUPLICATE_4dae_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_28_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_8fa7_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_29_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_b6d5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output, 32);
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_2_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l248_l244_l262_DUPLICATE_b3f8_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_30_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_6c97_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_31_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_b772_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_32_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_1a11_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_33_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_70f2_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_34_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_8029_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_35_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_bb47_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_36_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_4765_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_37_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_75bc_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_38_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_57c2_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_39_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_b3fb_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output, 32);
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_3_d41d_chacha20poly1305_decrypt_tb_c_l244_l234_l262_l248_l254_DUPLICATE_40ed_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_40_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l234_l262_DUPLICATE_e557_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_41_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_9498_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_42_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_6861_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_43_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_e107_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_44_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_4df3_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_45_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_1449_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_46_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_1c66_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_47_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2443_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_48_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_e555_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_49_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_caa5_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output, 32);
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_4_d41d_chacha20poly1305_decrypt_tb_c_l248_l234_l254_l244_l262_DUPLICATE_d04f_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_50_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_42c6_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_51_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_7e1c_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_52_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e10_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_53_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0849_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_54_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_7a4c_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_55_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0497_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_56_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_4323_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_57_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_e5c8_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_58_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_f737_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_59_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_2ff1_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output, 32);
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_5_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l234_l244_l254_DUPLICATE_1487_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_60_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_7c56_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_61_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_388a_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_62_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_16b9_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_63_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_617c_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_64_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_732a_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_65_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_eada_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_66_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_ceba_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_67_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_a55c_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_68_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_a5ec_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_69_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l254_l266_DUPLICATE_6aef_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output, 32);
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_6_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l234_l254_DUPLICATE_a270_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_70_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l254_l262_DUPLICATE_e1b4_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_71_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l266_l234_DUPLICATE_617e_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_72_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l266_l262_DUPLICATE_d93f_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_73_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_df0b_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_74_d41d_chacha20poly1305_decrypt_tb_c_l234_l262_l254_l266_DUPLICATE_a20d_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_75_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_9864_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_76_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_2818_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_77_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_4f4b_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_78_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l234_l262_DUPLICATE_d888_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_79_d41d_chacha20poly1305_decrypt_tb_c_l266_l254_l262_l234_DUPLICATE_2466_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output, 32);
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_7_d41d_chacha20poly1305_decrypt_tb_c_l234_l248_l254_l244_l262_DUPLICATE_6dbf_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_80_d41d_chacha20poly1305_decrypt_tb_c_l262_l254_l234_l266_DUPLICATE_77ac_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_81_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_0cc4_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_82_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_1da5_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_83_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_210e_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_84_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_51b7_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_85_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_9333_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_86_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_0ad3_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_87_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_2d4e_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_88_d41d_chacha20poly1305_decrypt_tb_c_l234_l254_l262_l266_DUPLICATE_3aa9_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_89_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l254_l234_DUPLICATE_f361_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output, 32);
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_8_d41d_chacha20poly1305_decrypt_tb_c_l244_l262_l248_l254_l234_DUPLICATE_c586_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_90_d41d_chacha20poly1305_decrypt_tb_c_l254_l262_l234_l266_DUPLICATE_5eb0_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_91_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_4d6c_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_92_d41d_chacha20poly1305_decrypt_tb_c_l266_l262_l234_l254_DUPLICATE_7a76_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_93_d41d_chacha20poly1305_decrypt_tb_c_l262_l234_l266_l254_DUPLICATE_b23f_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_94_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_42b2_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_95_d41d_chacha20poly1305_decrypt_tb_c_l266_l234_l262_l254_DUPLICATE_55f1_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_96_d41d_chacha20poly1305_decrypt_tb_c_l254_l234_l262_l266_DUPLICATE_5543_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_97_d41d_chacha20poly1305_decrypt_tb_c_l262_l266_l234_l254_DUPLICATE_4e14_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_98_d41d_chacha20poly1305_decrypt_tb_c_l234_l266_l262_l254_DUPLICATE_d818_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_99_d41d_chacha20poly1305_decrypt_tb_c_l254_l266_l262_l234_DUPLICATE_24aa_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right := VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 := resize(VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output, 32);
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse := VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue := VAR_CONST_REF_RD_char_char_128_9_d41d_chacha20poly1305_decrypt_tb_c_l248_l262_l244_l234_l254_DUPLICATE_7383_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_0_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l209_l220_DUPLICATE_114b_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_100_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_0841_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_101_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_948a_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_102_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_d1f0_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_103_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_2625_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_104_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_60e0_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_105_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_907f_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_106_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_41f5_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_107_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_1b22_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_108_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_baba_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_109_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_b585_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_10_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_5931_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_110_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_c801_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_111_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_c43c_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_112_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_3449_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_113_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_b2c7_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_114_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_706b_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_115_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_55d7_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_116_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_2843_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_117_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_5f73_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_118_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_399f_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_119_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_f076_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_11_d41d_chacha20poly1305_decrypt_tb_c_l209_l216_l200_l220_DUPLICATE_6b2f_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_120_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_793e_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_121_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l216_l200_DUPLICATE_5b24_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_122_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_5ee1_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_123_d41d_chacha20poly1305_decrypt_tb_c_l226_l220_l200_l216_DUPLICATE_6409_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_124_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_2726_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_125_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_53c1_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_126_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_f0c7_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_127_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_a367_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_12_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l209_l220_DUPLICATE_3c33_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_13_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l209_DUPLICATE_0a9c_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_14_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l209_DUPLICATE_e585_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_15_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_76c9_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_16_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_37b3_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_17_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_0131_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_18_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_b125_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_19_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_27ec_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_1_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l209_l200_DUPLICATE_ea2b_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_20_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_bad5_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_21_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_d34a_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_22_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_2893_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_23_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_d3d5_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_24_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_233d_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_25_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_ede1_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_26_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_6ca5_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_27_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_88d4_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_28_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_dcf2_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_29_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_6d1b_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_2_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l216_l220_DUPLICATE_05db_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_30_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_212e_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_31_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_81c2_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_32_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_274d_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_33_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_648f_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_34_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_d8d5_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_35_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_a2f5_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_36_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_9187_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_37_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_c31b_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_38_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_e743_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_39_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_1d93_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_3_d41d_chacha20poly1305_decrypt_tb_c_l200_l209_l220_l216_DUPLICATE_67d2_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_40_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_7d1b_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_41_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_a62b_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_42_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_0d29_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_43_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_eded_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_44_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_6921_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_45_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_2ebd_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_46_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_d638_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_47_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_3b2d_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_48_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_18f4_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_49_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_7905_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_4_d41d_chacha20poly1305_decrypt_tb_c_l216_l209_l220_l200_DUPLICATE_f98f_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_50_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_8bee_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_51_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_d73b_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_52_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_8dd6_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_53_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_344b_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_54_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_6ad5_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_55_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_45df_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_56_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_e58b_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_57_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l220_l216_DUPLICATE_623d_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_58_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_b31b_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_59_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_0b54_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_5_d41d_chacha20poly1305_decrypt_tb_c_l209_l220_l200_l216_DUPLICATE_0fa2_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_60_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l200_l220_DUPLICATE_661d_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_61_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_160f_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_62_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_9900_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_63_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_dc0d_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_64_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_041f_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_65_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l226_l200_DUPLICATE_c563_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_66_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l226_DUPLICATE_d7f9_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_67_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_2e8e_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_68_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_9b84_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_69_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_f2fc_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_6_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l209_DUPLICATE_c74c_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_70_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l226_l216_DUPLICATE_62c5_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_71_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_4eac_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_72_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_2681_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_73_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_c522_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_74_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l216_l226_DUPLICATE_ec33_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_75_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l216_l220_DUPLICATE_16ac_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_76_d41d_chacha20poly1305_decrypt_tb_c_l216_l220_l200_l226_DUPLICATE_d355_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_77_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l220_l200_DUPLICATE_ae0d_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_78_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_399d_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_79_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6167_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_7_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l220_l209_DUPLICATE_81f7_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_80_d41d_chacha20poly1305_decrypt_tb_c_l200_l220_l216_l226_DUPLICATE_891d_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_81_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_52a0_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_82_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l200_l226_DUPLICATE_3119_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_83_d41d_chacha20poly1305_decrypt_tb_c_l220_l200_l226_l216_DUPLICATE_30b2_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_84_d41d_chacha20poly1305_decrypt_tb_c_l200_l226_l216_l220_DUPLICATE_b3ae_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_85_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_d04e_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_86_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l200_l216_DUPLICATE_6f6a_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_87_d41d_chacha20poly1305_decrypt_tb_c_l220_l216_l226_l200_DUPLICATE_8fa2_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_88_d41d_chacha20poly1305_decrypt_tb_c_l226_l200_l220_l216_DUPLICATE_549c_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_89_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_cc26_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_8_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l209_DUPLICATE_9b25_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_90_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_3571_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_91_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_57e4_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_92_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_4da2_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_93_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l220_l226_DUPLICATE_ed58_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_94_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_79c4_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_95_d41d_chacha20poly1305_decrypt_tb_c_l200_l216_l226_l220_DUPLICATE_6b90_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_96_d41d_chacha20poly1305_decrypt_tb_c_l220_l226_l216_l200_DUPLICATE_ce53_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_97_d41d_chacha20poly1305_decrypt_tb_c_l226_l216_l200_l220_DUPLICATE_8e5e_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_98_d41d_chacha20poly1305_decrypt_tb_c_l216_l200_l226_l220_DUPLICATE_4a76_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_99_d41d_chacha20poly1305_decrypt_tb_c_l216_l226_l220_l200_DUPLICATE_49c1_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue := VAR_CONST_REF_RD_uint8_t_uint8_t_144_9_d41d_chacha20poly1305_decrypt_tb_c_l220_l209_l200_l216_DUPLICATE_32b2_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iftrue := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l261_c1_8ede_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l207_c16_98a8_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_112_CONST_REF_RD_uint8_t_uint8_t_144_128_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_113_CONST_REF_RD_uint8_t_uint8_t_144_129_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_114_CONST_REF_RD_uint8_t_uint8_t_144_130_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_115_CONST_REF_RD_uint8_t_uint8_t_144_131_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_116_CONST_REF_RD_uint8_t_uint8_t_144_132_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_117_CONST_REF_RD_uint8_t_uint8_t_144_133_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_118_CONST_REF_RD_uint8_t_uint8_t_144_134_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_119_CONST_REF_RD_uint8_t_uint8_t_144_135_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_120_CONST_REF_RD_uint8_t_uint8_t_144_136_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_121_CONST_REF_RD_uint8_t_uint8_t_144_137_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_122_CONST_REF_RD_uint8_t_uint8_t_144_138_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_123_CONST_REF_RD_uint8_t_uint8_t_144_139_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_124_CONST_REF_RD_uint8_t_uint8_t_144_140_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_125_CONST_REF_RD_uint8_t_uint8_t_144_141_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_126_CONST_REF_RD_uint8_t_uint8_t_144_142_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l226_c46_c57a_ITER_127_CONST_REF_RD_uint8_t_uint8_t_144_143_d41d_chacha20poly1305_decrypt_tb_c_l226_c173_b5dd_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l242_c16_321a_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_100_CONST_REF_RD_char_char_128_116_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_101_CONST_REF_RD_char_char_128_117_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_102_CONST_REF_RD_char_char_128_118_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_103_CONST_REF_RD_char_char_128_119_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_104_CONST_REF_RD_char_char_128_120_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_105_CONST_REF_RD_char_char_128_121_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_106_CONST_REF_RD_char_char_128_122_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_107_CONST_REF_RD_char_char_128_123_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_108_CONST_REF_RD_char_char_128_124_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_109_CONST_REF_RD_char_char_128_125_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_110_CONST_REF_RD_char_char_128_126_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_111_CONST_REF_RD_char_char_128_127_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_96_CONST_REF_RD_char_char_128_112_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_97_CONST_REF_RD_char_char_128_113_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_98_CONST_REF_RD_char_char_128_114_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse := VAR_FOR_chacha20poly1305_decrypt_tb_c_l266_c46_5d3f_ITER_99_CONST_REF_RD_char_char_128_115_d41d_chacha20poly1305_decrypt_tb_c_l266_c168_d9f8_return_output;
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l254_c1_0e8a_return_output;
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_right := VAR_UNARY_OP_NOT_chacha20poly1305_decrypt_tb_c_l272_c69_ec38_return_output;
     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l201_c1_1f18] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l262_c1_116d] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l255_c13_ead1] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l255_c1_a50b] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX[chacha20poly1305_decrypt_tb_c_l207_c13_1eb2] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output := FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l243_c1_fe25] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l257_c1_a633] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ[chacha20poly1305_decrypt_tb_c_l244_c20_3200] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l220_c13_2aef] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l262_c13_31d9] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS[chacha20poly1305_decrypt_tb_c_l246_c47_5882] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_left;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_right;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output;

     -- Submodule level 4
     VAR_printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l257_c1_a633_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_NEQ_chacha20poly1305_decrypt_tb_c_l244_c20_3200_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0 := resize(unsigned(std_logic_vector(VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_BIN_OP_PLUS_chacha20poly1305_decrypt_tb_c_l246_c47_5882_return_output)),32);
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l243_c1_fe25_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l201_c1_1f18_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l255_c1_a50b_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l262_c1_116d_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l220_c13_2aef_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l255_c13_ead1_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l262_c13_31d9_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_plaintext_pos_chacha20poly1305_decrypt_tb_c_l246_c30_af0f_0;
     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l217_c1_0485] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed[chacha20poly1305_decrypt_tb_c_l218_c62_4023] LATENCY=0
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l218_c62_4023_return_output := CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed(
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output);

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c(
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_0_chacha20poly1305_decrypt_axis_in_data_tdata_0_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_1_chacha20poly1305_decrypt_axis_in_data_tdata_1_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_2_chacha20poly1305_decrypt_axis_in_data_tdata_2_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_3_chacha20poly1305_decrypt_axis_in_data_tdata_3_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_4_chacha20poly1305_decrypt_axis_in_data_tdata_4_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_5_chacha20poly1305_decrypt_axis_in_data_tdata_5_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_6_chacha20poly1305_decrypt_axis_in_data_tdata_6_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_7_chacha20poly1305_decrypt_axis_in_data_tdata_7_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_8_chacha20poly1305_decrypt_axis_in_data_tdata_8_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_9_chacha20poly1305_decrypt_axis_in_data_tdata_9_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_10_chacha20poly1305_decrypt_axis_in_data_tdata_10_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_11_chacha20poly1305_decrypt_axis_in_data_tdata_11_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_12_chacha20poly1305_decrypt_axis_in_data_tdata_12_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_13_chacha20poly1305_decrypt_axis_in_data_tdata_13_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_14_chacha20poly1305_decrypt_axis_in_data_tdata_14_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     to_unsigned(1, 1),
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l203_c9_9137_ITER_15_chacha20poly1305_decrypt_axis_in_data_tdata_15_MUX_chacha20poly1305_decrypt_tb_c_l207_c13_1eb2_return_output,
     VAR_BIN_OP_LTE_chacha20poly1305_decrypt_tb_c_l213_c56_ca58_return_output,
     to_unsigned(1, 1));

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96[chacha20poly1305_decrypt_tb_c_l263_c18_9c96] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_chacha20poly1305_decrypt_tb_c_l263_c18_9c96_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8[chacha20poly1305_decrypt_tb_c_l256_c17_35f8] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_chacha20poly1305_decrypt_tb_c_l256_c17_35f8_CLOCK_ENABLE;
     -- Inputs
     -- Outputs

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c[chacha20poly1305_decrypt_tb_c_l258_c17_2a1c] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_chacha20poly1305_decrypt_tb_c_l258_c17_2a1c_arg0;
     -- Outputs

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l245_c1_df10] LATENCY=0
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_cond;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iftrue;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_iffalse;
     -- Outputs
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output := FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l254_c9_e02a] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l216_c9_bce0] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;

     -- Submodule level 5
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE := VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l245_c1_df10_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l217_c1_0485_return_output;
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_chacha20poly1305_decrypt_axis_in_TRUE_INPUT_MUX_CONST_REF_RD_axis128_t_stream_t_axis128_t_stream_t_0c8c_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l216_c9_bce0_return_output;
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l254_c9_e02a_return_output;
     -- plaintext_out_expected_42_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_111_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_33_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_57_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_51_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_27_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_13_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_25_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_71_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_14_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_78_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_43_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_35_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_31_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_2_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_5_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- plaintext_out_expected_87_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_76_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_12_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_47_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_86_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_121_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_31_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_72_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_98_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_8_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- chacha20poly1305_decrypt_axis_in_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_61_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_43_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_91_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_113_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_68_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_108_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_104_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_87_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_60_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_46_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_52_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_82_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_64_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_30_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_103_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_68_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_84_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_39_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_63_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_57_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_101_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_50_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_0_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_15_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_45_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_99_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_76_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_44_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_107_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_10_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_88_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_80_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_54_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_112_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_105_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_24_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_28_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_85_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_62_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_99_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_35_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_81_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_49_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_14_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_109_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_126_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_0_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_86_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_106_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_123_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_36_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_25_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_110_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_40_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_93_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_32_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_58_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_107_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_70_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_125_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_79_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_102_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_96_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_94_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_24_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_72_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_1_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_118_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_95_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_50_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_38_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_10_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_20_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_28_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_79_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_6_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_70_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_75_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_41_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_7_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_46_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_101_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_64_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_89_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_106_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_2_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_2_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_12_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_29_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_110_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_4_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_92_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_20_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_85_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_55_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_98_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_23_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_34_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_45_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_6_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- plaintext_out_expected_13_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_115_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_65_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_94_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_3_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- plaintext_out_expected_82_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_26_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_33_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_8_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_53_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_62_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_97_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_48_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_92_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_44_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_22_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_56_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_88_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- uint8_array16_be[chacha20poly1305_decrypt_tb_c_l218_c45_791a] LATENCY=0
     VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l218_c45_791a_return_output := uint8_array16_be(
     VAR_CONST_REF_RD_uint8_t_16_axis128_t_stream_t_data_tdata_deed_chacha20poly1305_decrypt_tb_c_l218_c62_4023_return_output);

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_7_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_103_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_66_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_29_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_15_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_73_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_90_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_0_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_100_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_56_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_11_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_54_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l220_c1_ea25] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output;

     -- ciphertext_in_stream_48_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_41_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_13_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_61_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_21_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_102_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- input_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_90_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_59_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_27_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_16_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_21_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_40_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_78_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_80_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_3_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_42_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_53_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_120_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_17_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_67_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_4_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_47_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_9_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_91_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_67_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_11_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- plaintext_out_expected_18_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_10_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- plaintext_out_expected_77_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_93_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_9_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_26_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_104_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_5_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_18_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_22_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_124_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_97_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_11_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_111_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_59_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_119_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_49_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_1_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_12_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_38_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_19_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_100_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_75_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_83_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_23_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_63_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_127_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_116_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_15_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_73_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_74_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_81_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_74_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_19_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_55_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_6_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_69_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_71_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_69_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_37_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_4_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- plaintext_out_expected_37_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_39_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_16_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_95_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_30_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_89_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_36_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_17_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_84_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_14_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_58_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_108_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_65_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_66_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_96_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951[chacha20poly1305_decrypt_tb_c_l247_c21_9951] LATENCY=0
     -- Clock enable
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_CLOCK_ENABLE;
     -- Inputs
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg0;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg1;
     FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2 <= VAR_FOR_chacha20poly1305_decrypt_tb_c_l240_c9_e2e7_ITER_9_printf_chacha20poly1305_decrypt_tb_c_l247_c21_9951_chacha20poly1305_decrypt_tb_c_l247_c21_9951_arg2;
     -- Outputs

     -- ciphertext_in_stream_83_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_105_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_3_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_7_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_32_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_77_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_60_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_122_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_5_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_52_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- ciphertext_in_stream_114_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_1_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_51_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_109_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- ciphertext_in_stream_117_MUX[chacha20poly1305_decrypt_tb_c_l200_c5_43ad] LATENCY=0
     -- Inputs
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_cond;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iftrue;
     ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse <= VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output := ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;

     -- plaintext_out_expected_34_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- plaintext_out_expected_8_MUX[chacha20poly1305_decrypt_tb_c_l234_c5_c0f6] LATENCY=0
     -- Inputs
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_cond;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iftrue;
     plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse <= VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output := plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;

     -- Submodule level 6
     VAR_printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l220_c1_ea25_return_output;
     REG_VAR_chacha20poly1305_decrypt_axis_in := VAR_chacha20poly1305_decrypt_axis_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_left := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_left := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_var_dim_0 := resize(VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output, 1);
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_var_dim_0 := resize(VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output, 1);
     REG_VAR_input_packet_count := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg0 := VAR_input_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output;
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_left := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output;
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l218_c45_791a_return_output;
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l218_c45_791a_return_output;
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l218_c45_791a_return_output;
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_x := VAR_uint8_array16_be_chacha20poly1305_decrypt_tb_c_l218_c45_791a_return_output;
     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l272_c9_d81d] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output;

     -- CONST_SR_32[chacha20poly1305_decrypt_tb_c_l218_c237_3380] LATENCY=0
     -- Inputs
     CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_x <= VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_x;
     -- Outputs
     VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output := CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output;

     -- CONST_SR_64[chacha20poly1305_decrypt_tb_c_l218_c207_36cf] LATENCY=0
     -- Inputs
     CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_x <= VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_x;
     -- Outputs
     VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output := CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output;

     -- VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8[chacha20poly1305_decrypt_tb_c_l289_c43_c7a8] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_0;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_1 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_ref_toks_1;
     VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_var_dim_0 <= VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output := VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output;

     -- CONST_REF_RD_uint8_t_144_uint8_t_144_10fa_chacha20poly1305_decrypt_tb_c_l286_l283_l272_DUPLICATE_f8a4 LATENCY=0
     VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_10fa_chacha20poly1305_decrypt_tb_c_l286_l283_l272_DUPLICATE_f8a4_return_output := CONST_REF_RD_uint8_t_144_uint8_t_144_10fa(
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
     VAR_ciphertext_in_stream_100_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_45_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_109_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_118_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_11_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_75_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_20_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_84_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_29_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_93_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_38_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_102_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_47_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_111_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_4_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_68_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_13_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_77_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_22_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_86_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_31_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_95_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_40_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_104_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_61_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_6_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_125_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_70_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_15_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_79_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_24_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_88_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_33_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_97_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_54_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_63_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_8_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_127_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_72_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_17_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_81_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_26_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_90_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_56_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_1_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_120_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_65_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_10_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_74_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_19_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_83_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_28_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_92_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_49_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_113_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_58_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_3_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_122_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_67_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_12_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_76_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_21_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_85_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_42_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_106_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_51_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_115_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_60_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_5_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_124_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_69_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_14_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_78_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_35_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_99_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_44_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_108_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_53_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_117_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_62_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_7_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_126_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_71_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_37_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_101_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_46_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_110_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_55_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_0_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_119_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_64_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_73_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_30_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_94_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_39_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_103_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_48_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_112_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_57_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_2_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_121_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_66_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_23_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_87_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_32_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_96_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_41_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_105_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_50_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_114_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_59_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_123_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_16_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_80_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_25_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_89_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_34_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_98_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_43_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_107_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_52_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_116_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_9_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_18_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_82_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_27_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_91_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output,
     VAR_ciphertext_in_stream_36_MUX_chacha20poly1305_decrypt_tb_c_l200_c5_43ad_return_output);

     -- CONST_SR_0[chacha20poly1305_decrypt_tb_c_l218_c267_24cf] LATENCY=0
     -- Inputs
     CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_x <= VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_x;
     -- Outputs
     VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output := CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0[chacha20poly1305_decrypt_tb_c_l221_c17_56b0] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_chacha20poly1305_decrypt_tb_c_l221_c17_56b0_arg0;
     -- Outputs

     -- CONST_REF_RD_char_128_char_128_1091_chacha20poly1305_decrypt_tb_c_l283_l272_l286_DUPLICATE_d4fa LATENCY=0
     VAR_CONST_REF_RD_char_128_char_128_1091_chacha20poly1305_decrypt_tb_c_l283_l272_l286_DUPLICATE_d4fa_return_output := CONST_REF_RD_char_128_char_128_1091(
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l173_c5_dd91_return_output,
     VAR_plaintext_out_expected_108_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_53_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_50_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_62_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_59_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_4_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_68_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_13_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_77_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_22_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_19_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_86_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_83_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_28_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_92_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_37_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_101_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_46_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_110_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_55_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_52_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_61_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_6_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_70_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_15_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_12_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_79_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_76_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_21_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_88_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_85_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_30_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_94_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_39_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_103_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_48_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_45_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_109_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_54_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_63_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_8_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_5_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_72_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_17_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_69_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_14_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_81_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_78_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_23_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_87_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_32_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_96_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_41_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_105_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_38_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_102_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_47_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_111_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_56_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_1_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_65_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_10_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_7_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_74_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_71_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_16_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_80_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_25_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_89_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_34_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_98_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_31_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_43_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_95_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_107_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_40_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_104_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_49_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_58_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_3_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_0_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_67_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_64_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_9_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_73_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_18_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_82_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_27_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_91_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_24_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_36_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_100_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_33_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_97_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_42_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_106_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_51_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_60_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_57_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_2_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_66_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_11_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_75_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_20_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_84_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_29_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_93_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_26_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_90_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_35_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_99_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output,
     VAR_plaintext_out_expected_44_MUX_chacha20poly1305_decrypt_tb_c_l234_c5_c0f6_return_output);

     -- VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8[chacha20poly1305_decrypt_tb_c_l288_c40_1f85] LATENCY=0
     -- Inputs
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_0;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_1 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_ref_toks_1;
     VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_var_dim_0 <= VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_var_dim_0;
     -- Outputs
     VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output := VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output;

     -- BIN_OP_EQ[chacha20poly1305_decrypt_tb_c_l286_c17_1b46] LATENCY=0
     -- Inputs
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_left <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_left;
     BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_right <= VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_right;
     -- Outputs
     VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output := BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;

     -- CONST_SR_96[chacha20poly1305_decrypt_tb_c_l218_c176_9ef3] LATENCY=0
     -- Inputs
     CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_x <= VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_x;
     -- Outputs
     VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output := CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output;

     -- Submodule level 7
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_left := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l272_c9_d81d_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond := VAR_BIN_OP_EQ_chacha20poly1305_decrypt_tb_c_l286_c17_1b46_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := VAR_CONST_REF_RD_char_128_char_128_1091_chacha20poly1305_decrypt_tb_c_l283_l272_l286_DUPLICATE_d4fa_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse := VAR_CONST_REF_RD_char_128_char_128_1091_chacha20poly1305_decrypt_tb_c_l283_l272_l286_DUPLICATE_d4fa_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse := VAR_CONST_REF_RD_char_128_char_128_1091_chacha20poly1305_decrypt_tb_c_l283_l272_l286_DUPLICATE_d4fa_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_10fa_chacha20poly1305_decrypt_tb_c_l286_l283_l272_DUPLICATE_f8a4_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_10fa_chacha20poly1305_decrypt_tb_c_l286_l283_l272_DUPLICATE_f8a4_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse := VAR_CONST_REF_RD_uint8_t_144_uint8_t_144_10fa_chacha20poly1305_decrypt_tb_c_l286_l283_l272_DUPLICATE_f8a4_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg3 := resize(VAR_CONST_SR_0_chacha20poly1305_decrypt_tb_c_l218_c267_24cf_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg2 := resize(VAR_CONST_SR_32_chacha20poly1305_decrypt_tb_c_l218_c237_3380_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg1 := resize(VAR_CONST_SR_64_chacha20poly1305_decrypt_tb_c_l218_c207_36cf_return_output, 32);
     VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg0 := resize(VAR_CONST_SR_96_chacha20poly1305_decrypt_tb_c_l218_c176_9ef3_return_output, 32);
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg1 := VAR_VAR_REF_RD_uint32_t_uint32_t_2_VAR_90b8_chacha20poly1305_decrypt_tb_c_l289_c43_c7a8_return_output;
     VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l288_c17_9f8c := VAR_VAR_REF_RD_uint8_t_144_uint8_t_2_144_VAR_90b8_chacha20poly1305_decrypt_tb_c_l288_c40_1f85_return_output.data;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue := VAR_ciphertext_in_stream_chacha20poly1305_decrypt_tb_c_l288_c17_9f8c;
     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l272_c9_c63b] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;

     -- printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25[chacha20poly1305_decrypt_tb_c_l218_c108_dc25] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg1;
     printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg2 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg2;
     printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg3 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_chacha20poly1305_decrypt_tb_c_l218_c108_dc25_arg3;
     -- Outputs

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l286_c13_9fea] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;

     -- Submodule level 8
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_left := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_c63b_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l286_c13_9fea_return_output;
     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;

     -- BIN_OP_AND[chacha20poly1305_decrypt_tb_c_l272_c9_dd50] LATENCY=0
     -- Inputs
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_left <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_left;
     BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_right <= VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_right;
     -- Outputs
     VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output := BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;

     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l283_c9_93c2] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;

     -- Submodule level 9
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond := VAR_BIN_OP_AND_chacha20poly1305_decrypt_tb_c_l272_c9_dd50_return_output;
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l283_c9_93c2_return_output;
     -- plaintext_out_size_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- plaintext_remaining_out_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- output_packet_count_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l273_c1_c4e6] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output;

     -- ciphertext_remaining_in_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- plaintext_out_expected_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- ciphertext_in_stream_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l272_c5_0dda] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;

     -- Submodule level 10
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iffalse := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l273_c1_c4e6_return_output;
     REG_VAR_ciphertext_in_stream := VAR_ciphertext_in_stream_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     REG_VAR_ciphertext_remaining_in := VAR_ciphertext_remaining_in_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_right := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     REG_VAR_output_packet_count := VAR_output_packet_count_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     REG_VAR_plaintext_out_expected := VAR_plaintext_out_expected_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     REG_VAR_plaintext_out_size := VAR_plaintext_out_size_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     REG_VAR_plaintext_remaining_out := VAR_plaintext_remaining_out_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iffalse := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l272_c5_0dda_return_output;
     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l275_c1_e50f] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output;

     -- BIN_OP_GT[chacha20poly1305_decrypt_tb_c_l305_c9_276d] LATENCY=0
     -- Inputs
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_left <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_left;
     BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_right <= VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_right;
     -- Outputs
     VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output := BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output;

     -- FALSE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l277_c1_ea4e] LATENCY=0
     -- Inputs
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_cond <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_cond;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iftrue <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iftrue;
     FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iffalse <= VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_iffalse;
     -- Outputs
     VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output := FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output;

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l284_c1_88f0] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output;

     -- Submodule level 11
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_cond := VAR_BIN_OP_GT_chacha20poly1305_decrypt_tb_c_l305_c9_276d_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_CLOCK_ENABLE := VAR_FALSE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l277_c1_ea4e_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l275_c1_e50f_return_output;
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iftrue := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l284_c1_88f0_return_output;
     -- printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7[chacha20poly1305_decrypt_tb_c_l276_c13_2af7] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_chacha20poly1305_decrypt_tb_c_l276_c13_2af7_arg0;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87[chacha20poly1305_decrypt_tb_c_l278_c13_ab87] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_chacha20poly1305_decrypt_tb_c_l278_c13_ab87_arg0;
     -- Outputs

     -- TRUE_CLOCK_ENABLE_MUX[chacha20poly1305_decrypt_tb_c_l286_c1_c205] LATENCY=0
     -- Inputs
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_cond <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_cond;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iftrue <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iftrue;
     TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iffalse <= VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_iffalse;
     -- Outputs
     VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output := TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output;

     -- tag_match_checked_MUX[chacha20poly1305_decrypt_tb_c_l305_c5_427d] LATENCY=0
     -- Inputs
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_cond <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_cond;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iftrue <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iftrue;
     tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iffalse <= VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_iffalse;
     -- Outputs
     VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output := tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output;

     -- Submodule level 12
     VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output;
     VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_CLOCK_ENABLE := VAR_TRUE_CLOCK_ENABLE_MUX_chacha20poly1305_decrypt_tb_c_l286_c1_c205_return_output;
     REG_VAR_tag_match_checked := VAR_tag_match_checked_MUX_chacha20poly1305_decrypt_tb_c_l305_c5_427d_return_output;
     -- printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9[chacha20poly1305_decrypt_tb_c_l298_c17_cae9] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_chacha20poly1305_decrypt_tb_c_l298_c17_cae9_arg1;
     -- Outputs

     -- printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec[chacha20poly1305_decrypt_tb_c_l290_c17_c7ec] LATENCY=0
     -- Clock enable
     printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_CLOCK_ENABLE <= VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_CLOCK_ENABLE;
     -- Inputs
     printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg0 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg0;
     printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg1 <= VAR_printf_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_chacha20poly1305_decrypt_tb_c_l290_c17_c7ec_arg1;
     -- Outputs

     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

-- Write regs vars to comb logic
REG_COMB_input_packet_count <= REG_VAR_input_packet_count;
REG_COMB_ciphertext_in_stream <= REG_VAR_ciphertext_in_stream;
REG_COMB_ciphertext_remaining_in <= REG_VAR_ciphertext_remaining_in;
REG_COMB_cycle_counter <= REG_VAR_cycle_counter;
REG_COMB_output_packet_count <= REG_VAR_output_packet_count;
REG_COMB_plaintext_out_size <= REG_VAR_plaintext_out_size;
REG_COMB_plaintext_remaining_out <= REG_VAR_plaintext_remaining_out;
REG_COMB_plaintext_out_expected <= REG_VAR_plaintext_out_expected;
REG_COMB_tag_match_checked <= REG_VAR_tag_match_checked;
REG_COMB_chacha20poly1305_decrypt_axis_in <= REG_VAR_chacha20poly1305_decrypt_axis_in;
-- Global wires driven various places in pipeline
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_key <= VAR_chacha20poly1305_decrypt_key;
else
  module_to_global.chacha20poly1305_decrypt_key <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_nonce <= VAR_chacha20poly1305_decrypt_nonce;
else
  module_to_global.chacha20poly1305_decrypt_nonce <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad <= VAR_chacha20poly1305_decrypt_aad;
else
  module_to_global.chacha20poly1305_decrypt_aad <= (others => to_unsigned(0, 8));
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_aad_len <= VAR_chacha20poly1305_decrypt_aad_len;
else
  module_to_global.chacha20poly1305_decrypt_aad_len <= to_unsigned(0, 8);
end if;
if clk_en_internal='1' then
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= VAR_chacha20poly1305_decrypt_axis_out_ready;
else
  module_to_global.chacha20poly1305_decrypt_axis_out_ready <= to_unsigned(0, 1);
end if;
end process;

-- Register comb signals
process(clk) is
begin
 if rising_edge(clk) then
 if clk_en_internal='1' then
     input_packet_count <= REG_COMB_input_packet_count;
     ciphertext_in_stream <= REG_COMB_ciphertext_in_stream;
     ciphertext_remaining_in <= REG_COMB_ciphertext_remaining_in;
     cycle_counter <= REG_COMB_cycle_counter;
     output_packet_count <= REG_COMB_output_packet_count;
     plaintext_out_size <= REG_COMB_plaintext_out_size;
     plaintext_remaining_out <= REG_COMB_plaintext_remaining_out;
     plaintext_out_expected <= REG_COMB_plaintext_out_expected;
     tag_match_checked <= REG_COMB_tag_match_checked;
     chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in;
 end if;
 end if;
end process;
-- Shared global regs
module_to_global.chacha20poly1305_decrypt_axis_in <= REG_COMB_chacha20poly1305_decrypt_axis_in when clk_en_internal='1' else chacha20poly1305_decrypt_axis_in;

end arch;
