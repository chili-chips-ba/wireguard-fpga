-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 16
entity axis128_keep_count_0CLK_08de2a73 is
port(
 axis : in axis128_t;
 return_output : out unsigned(4 downto 0));
end axis128_keep_count_0CLK_08de2a73;
architecture arch of axis128_keep_count_0CLK_08de2a73 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_2c77]
signal FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_efc2]
signal FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_c9fe]
signal FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_7e8f]
signal FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_5c59]
signal FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_7411]
signal FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_e7eb]
signal FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_c9b6]
signal FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_5cd8]
signal FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_3e67]
signal FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_47f1]
signal FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_e153]
signal FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_94e9]
signal FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_82fe]
signal FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_0844]
signal FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output : unsigned(5 downto 0);

-- FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_cc71]
signal FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_left : unsigned(4 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_right : unsigned(0 downto 0);
signal FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output : unsigned(5 downto 0);


begin

-- SUBMODULE INSTANCES 
-- FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_left,
FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_right,
FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_left,
FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_right,
FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_left,
FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_right,
FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_left,
FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_right,
FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_left,
FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_right,
FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_left,
FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_right,
FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_left,
FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_right,
FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_left,
FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_right,
FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_left,
FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_right,
FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_left,
FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_right,
FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_left,
FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_right,
FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_left,
FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_right,
FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_left,
FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_right,
FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_left,
FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_right,
FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_left,
FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_right,
FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output);

-- FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71 : 0 clocks latency
FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71 : entity work.BIN_OP_PLUS_uint5_t_uint1_t_0CLK_de264c78 port map (
FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_left,
FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_right,
FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 axis,
 -- All submodule outputs
 FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output,
 FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output,
 FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output,
 FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output,
 FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output,
 FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output,
 FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output,
 FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output,
 FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output,
 FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output,
 FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output,
 FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output,
 FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output,
 FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output,
 FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output,
 FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(4 downto 0);
 variable VAR_axis : axis128_t;
 variable VAR_rv : unsigned(4 downto 0);
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_0_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_1_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_2_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_3_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_4_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_5_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_6_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_7_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_8_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_9_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_10_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_11_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_12_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_13_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_14_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output : unsigned(5 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_15_rv_axis_h_l91_c5_dd39 : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_left : unsigned(4 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_11b5_return_output : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_right : unsigned(0 downto 0);
 variable VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output : unsigned(5 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_left := to_unsigned(0, 5);

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_axis := axis;

     -- Submodule level 0
     -- FOR_axis_h_l90_c3_7193_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(4);

     -- FOR_axis_h_l90_c3_7193_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(5);

     -- FOR_axis_h_l90_c3_7193_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(14);

     -- FOR_axis_h_l90_c3_7193_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(2);

     -- FOR_axis_h_l90_c3_7193_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(1);

     -- FOR_axis_h_l90_c3_7193_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(11);

     -- FOR_axis_h_l90_c3_7193_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(6);

     -- FOR_axis_h_l90_c3_7193_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(10);

     -- FOR_axis_h_l90_c3_7193_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(0);

     -- FOR_axis_h_l90_c3_7193_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(9);

     -- FOR_axis_h_l90_c3_7193_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(8);

     -- FOR_axis_h_l90_c3_7193_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(15);

     -- FOR_axis_h_l90_c3_7193_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(13);

     -- FOR_axis_h_l90_c3_7193_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(7);

     -- FOR_axis_h_l90_c3_7193_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(3);

     -- FOR_axis_h_l90_c3_7193_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d[axis_h_l91_c11_11b5] LATENCY=0
     VAR_FOR_axis_h_l90_c3_7193_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_11b5_return_output := VAR_axis.tkeep(12);

     -- Submodule level 1
     VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_right := VAR_FOR_axis_h_l90_c3_7193_ITER_0_CONST_REF_RD_uint1_t_axis128_t_tkeep_0_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_right := VAR_FOR_axis_h_l90_c3_7193_ITER_10_CONST_REF_RD_uint1_t_axis128_t_tkeep_10_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_right := VAR_FOR_axis_h_l90_c3_7193_ITER_11_CONST_REF_RD_uint1_t_axis128_t_tkeep_11_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_right := VAR_FOR_axis_h_l90_c3_7193_ITER_12_CONST_REF_RD_uint1_t_axis128_t_tkeep_12_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_right := VAR_FOR_axis_h_l90_c3_7193_ITER_13_CONST_REF_RD_uint1_t_axis128_t_tkeep_13_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_right := VAR_FOR_axis_h_l90_c3_7193_ITER_14_CONST_REF_RD_uint1_t_axis128_t_tkeep_14_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_right := VAR_FOR_axis_h_l90_c3_7193_ITER_15_CONST_REF_RD_uint1_t_axis128_t_tkeep_15_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_right := VAR_FOR_axis_h_l90_c3_7193_ITER_1_CONST_REF_RD_uint1_t_axis128_t_tkeep_1_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_right := VAR_FOR_axis_h_l90_c3_7193_ITER_2_CONST_REF_RD_uint1_t_axis128_t_tkeep_2_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_right := VAR_FOR_axis_h_l90_c3_7193_ITER_3_CONST_REF_RD_uint1_t_axis128_t_tkeep_3_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_right := VAR_FOR_axis_h_l90_c3_7193_ITER_4_CONST_REF_RD_uint1_t_axis128_t_tkeep_4_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_right := VAR_FOR_axis_h_l90_c3_7193_ITER_5_CONST_REF_RD_uint1_t_axis128_t_tkeep_5_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_right := VAR_FOR_axis_h_l90_c3_7193_ITER_6_CONST_REF_RD_uint1_t_axis128_t_tkeep_6_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_right := VAR_FOR_axis_h_l90_c3_7193_ITER_7_CONST_REF_RD_uint1_t_axis128_t_tkeep_7_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_right := VAR_FOR_axis_h_l90_c3_7193_ITER_8_CONST_REF_RD_uint1_t_axis128_t_tkeep_8_d41d_axis_h_l91_c11_11b5_return_output;
     VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_right := VAR_FOR_axis_h_l90_c3_7193_ITER_9_CONST_REF_RD_uint1_t_axis128_t_tkeep_9_d41d_axis_h_l91_c11_11b5_return_output;
     -- FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS[axis_h_l91_c5_2c77] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_left;
     FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output := FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output;

     -- Submodule level 2
     VAR_FOR_axis_h_l90_c3_7193_ITER_0_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_0_BIN_OP_PLUS_axis_h_l91_c5_2c77_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_left := VAR_FOR_axis_h_l90_c3_7193_ITER_0_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS[axis_h_l91_c5_efc2] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_left;
     FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output := FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output;

     -- Submodule level 3
     VAR_FOR_axis_h_l90_c3_7193_ITER_1_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_1_BIN_OP_PLUS_axis_h_l91_c5_efc2_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_left := VAR_FOR_axis_h_l90_c3_7193_ITER_1_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS[axis_h_l91_c5_c9fe] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_left;
     FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output := FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output;

     -- Submodule level 4
     VAR_FOR_axis_h_l90_c3_7193_ITER_2_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_2_BIN_OP_PLUS_axis_h_l91_c5_c9fe_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_left := VAR_FOR_axis_h_l90_c3_7193_ITER_2_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS[axis_h_l91_c5_7e8f] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_left;
     FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output := FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output;

     -- Submodule level 5
     VAR_FOR_axis_h_l90_c3_7193_ITER_3_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_3_BIN_OP_PLUS_axis_h_l91_c5_7e8f_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_left := VAR_FOR_axis_h_l90_c3_7193_ITER_3_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS[axis_h_l91_c5_5c59] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_left;
     FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output := FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output;

     -- Submodule level 6
     VAR_FOR_axis_h_l90_c3_7193_ITER_4_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_4_BIN_OP_PLUS_axis_h_l91_c5_5c59_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_left := VAR_FOR_axis_h_l90_c3_7193_ITER_4_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS[axis_h_l91_c5_7411] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_left;
     FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output := FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output;

     -- Submodule level 7
     VAR_FOR_axis_h_l90_c3_7193_ITER_5_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_5_BIN_OP_PLUS_axis_h_l91_c5_7411_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_left := VAR_FOR_axis_h_l90_c3_7193_ITER_5_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS[axis_h_l91_c5_e7eb] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_left;
     FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output := FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output;

     -- Submodule level 8
     VAR_FOR_axis_h_l90_c3_7193_ITER_6_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_6_BIN_OP_PLUS_axis_h_l91_c5_e7eb_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_left := VAR_FOR_axis_h_l90_c3_7193_ITER_6_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS[axis_h_l91_c5_c9b6] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_left;
     FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output := FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output;

     -- Submodule level 9
     VAR_FOR_axis_h_l90_c3_7193_ITER_7_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_7_BIN_OP_PLUS_axis_h_l91_c5_c9b6_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_left := VAR_FOR_axis_h_l90_c3_7193_ITER_7_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS[axis_h_l91_c5_5cd8] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_left;
     FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output := FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output;

     -- Submodule level 10
     VAR_FOR_axis_h_l90_c3_7193_ITER_8_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_8_BIN_OP_PLUS_axis_h_l91_c5_5cd8_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_left := VAR_FOR_axis_h_l90_c3_7193_ITER_8_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS[axis_h_l91_c5_3e67] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_left;
     FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output := FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output;

     -- Submodule level 11
     VAR_FOR_axis_h_l90_c3_7193_ITER_9_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_9_BIN_OP_PLUS_axis_h_l91_c5_3e67_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_left := VAR_FOR_axis_h_l90_c3_7193_ITER_9_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS[axis_h_l91_c5_47f1] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_left;
     FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output := FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output;

     -- Submodule level 12
     VAR_FOR_axis_h_l90_c3_7193_ITER_10_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_10_BIN_OP_PLUS_axis_h_l91_c5_47f1_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_left := VAR_FOR_axis_h_l90_c3_7193_ITER_10_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS[axis_h_l91_c5_e153] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_left;
     FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output := FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output;

     -- Submodule level 13
     VAR_FOR_axis_h_l90_c3_7193_ITER_11_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_11_BIN_OP_PLUS_axis_h_l91_c5_e153_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_left := VAR_FOR_axis_h_l90_c3_7193_ITER_11_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS[axis_h_l91_c5_94e9] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_left;
     FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output := FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output;

     -- Submodule level 14
     VAR_FOR_axis_h_l90_c3_7193_ITER_12_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_12_BIN_OP_PLUS_axis_h_l91_c5_94e9_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_left := VAR_FOR_axis_h_l90_c3_7193_ITER_12_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS[axis_h_l91_c5_82fe] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_left;
     FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output := FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output;

     -- Submodule level 15
     VAR_FOR_axis_h_l90_c3_7193_ITER_13_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_13_BIN_OP_PLUS_axis_h_l91_c5_82fe_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_left := VAR_FOR_axis_h_l90_c3_7193_ITER_13_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS[axis_h_l91_c5_0844] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_left;
     FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output := FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output;

     -- Submodule level 16
     VAR_FOR_axis_h_l90_c3_7193_ITER_14_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_14_BIN_OP_PLUS_axis_h_l91_c5_0844_return_output, 5);
     VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_left := VAR_FOR_axis_h_l90_c3_7193_ITER_14_rv_axis_h_l91_c5_dd39;
     -- FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS[axis_h_l91_c5_cc71] LATENCY=0
     -- Inputs
     FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_left <= VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_left;
     FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_right <= VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_right;
     -- Outputs
     VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output := FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output;

     -- Submodule level 17
     VAR_FOR_axis_h_l90_c3_7193_ITER_15_rv_axis_h_l91_c5_dd39 := resize(VAR_FOR_axis_h_l90_c3_7193_ITER_15_BIN_OP_PLUS_axis_h_l91_c5_cc71_return_output, 5);
     VAR_return_output := VAR_FOR_axis_h_l90_c3_7193_ITER_15_rv_axis_h_l91_c5_dd39;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
