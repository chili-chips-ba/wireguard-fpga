-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 96
entity uint320_mul_0CLK_babc4282 is
port(
 a : in u320_t;
 b : in u320_t;
 return_output : out u320_t);
end uint320_mul_0CLK_babc4282;
architecture arch of uint320_mul_0CLK_babc4282 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_c7dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_c6ec]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_56cc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_c3d3]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_4dd8]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_1713]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_03e8]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_4c26]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_4c03]
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_57a2]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_13fd]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_2f4e]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_edbc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_07ed]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_a961]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_e943]
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_e468]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_eb04]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_8177]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_dd7e]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_c2cd]
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_bec3]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_9f23]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_right : unsigned(0 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_d9c3]
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc]
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c]
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);

-- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_6597]
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_left : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_right : unsigned(63 downto 0);
signal FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output : unsigned(64 downto 0);

function CONST_REF_RD_u320_t_u320_t_4216( ref_toks_0 : unsigned;
 ref_toks_1 : unsigned;
 ref_toks_2 : unsigned;
 ref_toks_3 : unsigned;
 ref_toks_4 : unsigned) return u320_t is
 
  variable base : u320_t; 
  variable return_output : u320_t;
begin
      base.limbs(0) := ref_toks_0;
      base.limbs(1) := ref_toks_1;
      base.limbs(2) := ref_toks_2;
      base.limbs(3) := ref_toks_3;
      base.limbs(4) := ref_toks_4;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_left,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_right,
FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_left,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_right,
FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_left,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_right,
FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806 : entity work.MUX_uint1_t_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf : entity work.BIN_OP_LT_uint64_t_uint64_t_0CLK_380ecc95 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb : entity work.MUX_uint1_t_uint1_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23 : entity work.BIN_OP_PLUS_uint64_t_uint1_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_left,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_right,
FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc : entity work.BIN_OP_INFERRED_MULT_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left,
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right,
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left,
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right,
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output);

-- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597 : 0 clocks latency
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597 : entity work.BIN_OP_PLUS_uint64_t_uint64_t_0CLK_de264c78 port map (
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_left,
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_right,
FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 a,
 b,
 -- All submodule outputs
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output,
 FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : u320_t;
 variable VAR_a : u320_t;
 variable VAR_b : u320_t;
 variable VAR_temp : u320_t;
 variable VAR_i : signed(31 downto 0);
 variable VAR_carry : unsigned(63 downto 0);
 variable VAR_j : signed(31 downto 0);
 variable VAR_high : unsigned(63 downto 0);
 variable VAR_low : unsigned(63 downto 0);
 variable VAR_product : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_old_value : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_52bb_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_52bb_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_52bb_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_52bb_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_00fb_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_52bb_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_right : unsigned(0 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_c892_return_output : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output : unsigned(127 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output : unsigned(64 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_left : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_right : unsigned(63 downto 0);
 variable VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output : unsigned(64 downto 0);
 variable VAR_res : u320_t;
 variable VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_39b1_return_output : u320_t;
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_9b0b_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_014e_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_d022_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_c892_DUPLICATE_120c_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_c892_DUPLICATE_8299_return_output : unsigned(63 downto 0);
 variable VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e020_return_output : unsigned(63 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_right := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse := to_unsigned(0, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse := to_unsigned(0, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue := to_unsigned(1, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue := to_unsigned(1, 1);
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l128_c34_52bb] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_52bb_return_output := u320_t_NULL.limbs(4);

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l128_c34_52bb] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_52bb_return_output := u320_t_NULL.limbs(0);

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l128_c34_52bb] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_52bb_return_output := u320_t_NULL.limbs(1);

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l128_c34_52bb] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_52bb_return_output := u320_t_NULL.limbs(3);

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l128_c34_52bb] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_52bb_return_output := u320_t_NULL.limbs(2);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l128_c34_52bb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l128_c34_52bb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l128_c34_52bb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l128_c34_52bb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l128_c34_52bb_return_output;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_a := a;
     VAR_b := b;

     -- Submodule level 0
     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c45_00fb]_DUPLICATE_9b0b LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_9b0b_return_output := VAR_b.limbs(1);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c32_c892]_DUPLICATE_e020 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e020_return_output := VAR_a.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d[poly1305_h_l127_c45_00fb]_DUPLICATE_d022 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_d022_return_output := VAR_b.limbs(3);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c32_c892]_DUPLICATE_e36b LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output := VAR_a.limbs(0);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c45_00fb]_DUPLICATE_014e LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_014e_return_output := VAR_b.limbs(2);

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c45_00fb] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_00fb_return_output := VAR_b.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d[poly1305_h_l127_c32_c892]_DUPLICATE_8299 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_c892_DUPLICATE_8299_return_output := VAR_a.limbs(2);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d[poly1305_h_l127_c32_c892]_DUPLICATE_120c LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_c892_DUPLICATE_120c_return_output := VAR_a.limbs(1);

     -- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d[poly1305_h_l127_c32_c892] LATENCY=0
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_c892_return_output := VAR_a.limbs(4);

     -- CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d[poly1305_h_l127_c45_00fb]_DUPLICATE_49e8 LATENCY=0
     VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output := VAR_b.limbs(0);

     -- Submodule level 1
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e36b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_0_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_49e8_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_c892_DUPLICATE_120c_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_c892_DUPLICATE_120c_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_c892_DUPLICATE_120c_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c32_c892_DUPLICATE_120c_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_9b0b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_9b0b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_9b0b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_1_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_9b0b_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_c892_DUPLICATE_8299_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_c892_DUPLICATE_8299_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c32_c892_DUPLICATE_8299_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_014e_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_014e_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_2_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_014e_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e020_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c32_c892_DUPLICATE_e020_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_d022_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_CONST_REF_RD_uint64_t_u320_t_limbs_3_d41d_poly1305_h_l127_c45_00fb_DUPLICATE_d022_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c45_00fb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_CONST_REF_RD_uint64_t_u320_t_limbs_4_d41d_poly1305_h_l127_c32_c892_return_output;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT[poly1305_h_l127_c32_b9dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output;

     -- Submodule level 2
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_INFERRED_MULT_poly1305_h_l127_c32_b9dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_product_poly1305_h_l127_c22_5f93_0;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_product_poly1305_h_l127_c22_5f93_0;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- Submodule level 3
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_c7dc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- Submodule level 4
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_c7dc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;

     -- Submodule level 5
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l132_c21_c806_return_output;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- Submodule level 6
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_c6ec] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output;

     -- Submodule level 7
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_c6ec_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_56cc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output;

     -- Submodule level 8
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_56cc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- Submodule level 9
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_57a2] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output;

     -- Submodule level 10
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_57a2_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_c3d3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;

     -- Submodule level 11
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_c3d3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_4dd8] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output;

     -- Submodule level 12
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_4dd8_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_13fd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- Submodule level 13
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_13fd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_2f4e] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- Submodule level 14
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_2f4e_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_1713] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output;

     -- Submodule level 15
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_1713_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_e468] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_03e8] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- Submodule level 16
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_03e8_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_e468_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_edbc] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- Submodule level 17
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_edbc_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_07ed] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output;

     -- Submodule level 18
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_07ed_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_eb04] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l134_c13_4c26] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- Submodule level 19
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l134_c13_4c26_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_eb04_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_3_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_8177] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS[poly1305_h_l133_c13_4c03] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- Submodule level 20
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_BIN_OP_PLUS_poly1305_h_l133_c13_4c03_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_8177_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_4_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l134_c13_a961] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- Submodule level 21
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l134_c13_a961_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_2_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l132_c21_a4cf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_bec3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS[poly1305_h_l133_c13_e943] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output;

     -- Submodule level 22
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_BIN_OP_PLUS_poly1305_h_l133_c13_e943_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l132_c21_a4cf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_bec3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_3_low_poly1305_h_l133_c13_3abd;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l134_c13_dd7e] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l132_c21_c806] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT[poly1305_h_l134_c22_8abf] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;

     -- Submodule level 23
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l134_c13_dd7e_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_LT_poly1305_h_l134_c22_8abf_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l132_c21_c806_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_1_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX[poly1305_h_l134_c22_e0eb] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_cond;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iftrue;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_iffalse;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS[poly1305_h_l133_c13_c2cd] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output;

     -- Submodule level 24
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_BIN_OP_PLUS_poly1305_h_l133_c13_c2cd_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_MUX_poly1305_h_l134_c22_e0eb_return_output;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_2_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l134_c13_9f23] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output;

     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- Submodule level 25
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l134_c13_9f23_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_high_poly1305_h_l134_c13_6ee4;
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS[poly1305_h_l133_c13_d9c3] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output;

     -- Submodule level 26
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_BIN_OP_PLUS_poly1305_h_l133_c13_d9c3_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_1_low_poly1305_h_l133_c13_3abd;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l131_c19_b86c] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output;

     -- Submodule level 27
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17 := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l131_c19_b86c_return_output, 64);
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_left := VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l131_c13_8a17;
     -- FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS[poly1305_h_l133_c13_6597] LATENCY=0
     -- Inputs
     FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_left <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_left;
     FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_right <= VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_right;
     -- Outputs
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output := FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output;

     -- Submodule level 28
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd := resize(VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_BIN_OP_PLUS_poly1305_h_l133_c13_6597_return_output, 64);
     -- CONST_REF_RD_u320_t_u320_t_4216[poly1305_h_l141_c18_39b1] LATENCY=0
     VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_39b1_return_output := CONST_REF_RD_u320_t_u320_t_4216(
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_0_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd,
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_1_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd,
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_2_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd,
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_3_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd,
     VAR_FOR_poly1305_h_l120_c5_fe90_ITER_4_FOR_poly1305_h_l123_c9_8444_ITER_0_low_poly1305_h_l133_c13_3abd);

     -- Submodule level 29
     VAR_return_output := VAR_CONST_REF_RD_u320_t_u320_t_4216_poly1305_h_l141_c18_39b1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
